`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Technische Universität München (TUM) / Fraunhofer Institute for Applied and Integrated Security (AISEC)
// Engineer: Tobias Stelzer
// 
// Create Date: 06/14/2022 12:27:48 PM
// Design Name: PQ_OTBN
// Module Name: tb_otbn
// Project Name: 2022-MA-PQ-ALU-OpenTitan
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_otbn
    import prim_alert_pkg::*;
    import otbn_pkg::*;
    import otbn_reg_pkg::*;
    import tb_tl_ul_pkg::*;
    (
    
    );
    
// Parameter
    localparam bit                   Stub         = 1'b0;
    localparam regfile_e             RegFile      = RegFileFF;
    localparam logic [NumAlerts-1:0] AlertAsyncOn = {NumAlerts{1'b0}};
    
    // Default seed and permutation for URND LFSR
    localparam urnd_lfsr_seed_t       RndCnstUrndLfsrSeed      = RndCnstUrndLfsrSeedDefault;
    localparam urnd_chunk_lfsr_perm_t RndCnstUrndChunkLfsrPerm = RndCnstUrndChunkLfsrPermDefault;  
     
    localparam string                 log_path = "/home/t_stelzer/projects/aisec/opentitan/hw/vendor/aisec_otbn_pq/dv/sv/log/";
    localparam string                 mem_path = "/home/t_stelzer/projects/aisec/opentitan/hw/vendor/aisec_otbn_pq/dv/sv/";
    
    // Filehandle, clock cycle counter, readback data variable, teststate
    integer                                     f;   
    integer                                     cc;
    integer                                     cc_start;
    integer                                     cc_stop;
    integer                                     cc_count_dilithium;
    integer                                     cc_count_kyber;
    
    integer                                     cc_count_dilithium_indirect;
    integer                                     cc_count_kyber_indirect;
    
    integer                                     cc_count_dilithium_inv;
    integer                                     cc_count_kyber_inv;    
    
    integer                                     cc_count_dilithium_inv_indirect;
    integer                                     cc_count_kyber_inv_indirect;    
 
    integer                                     cc_count_falcon512_indirect;
    integer                                     cc_count_falcon1024_indirect;

    integer                                     cc_count_falcon512_inv_indirect;
    integer                                     cc_count_falcon1024_inv_indirect;

    integer                                     cc_count_dilithium_pointwise_mul;
    integer                                     cc_count_kyber_base_mul;
    integer                                     cc_count_falcon512_pointwise_mul;
    integer                                     cc_count_falcon1024_pointwise_mul;

    
    logic                       [31:0]          rdbk;
    string                                      teststate;  
    integer                                     error_count;
    
    // Clock and Reset
    logic                                       clk_i;
    logic                                       rst_ni;

    // Bus Signals    
    tlul_pkg::tl_h2d_t                          tl_i_d,tl_i_q;
    tlul_pkg::tl_d2h_t                          tl_o;
    logic                                       err_tl;
       
    // Inter-module signals
    logic                                       idle_o;
    
    // Interrupts
    logic                                       intr_done_o;
    
    // Alerts
    prim_alert_pkg::alert_rx_t [NumAlerts-1:0] alert_rx_i;
    prim_alert_pkg::alert_tx_t [NumAlerts-1:0] alert_tx_o;
    
    // Memory configuration
    prim_ram_1p_pkg::ram_1p_cfg_t ram_cfg_i;

    
    // EDN clock and interface
    logic                                       clk_edn_i;
    logic                                       rst_edn_ni;
    
    edn_pkg::edn_req_t                          edn_rnd_o;
    edn_pkg::edn_rsp_t                          edn_rnd_i;
    
    edn_pkg::edn_req_t                          edn_urnd_o;
    edn_pkg::edn_rsp_t                          edn_urnd_i;
    
   
    
    
    // DUT   
    otbn #(.Stub(Stub),
        .RegFile(RegFile),
        .AlertAsyncOn(AlertAsyncOn),
        
        // Default seed and permutation for URND LFSR
        .RndCnstUrndLfsrSeed(RndCnstUrndLfsrSeed),
        .RndCnstUrndChunkLfsrPerm(RndCnstUrndChunkLfsrPerm))
    DUT (
        .clk_i(clk_i),
        .rst_ni(rst_ni),
        
        .tl_i(tl_i_q),
        .tl_o(tl_o),
        
          // Inter-module signals
        .idle_o(idle_o),
        
          // Interrupts
        .intr_done_o(intr_done_o),
        
          // Alerts
        .alert_rx_i(alert_rx_i),
        .alert_tx_o(alert_tx_o),
        
          // Memory configuration
        .ram_cfg_i(ram_cfg_i),
        
          // EDN clock and interface
        .clk_edn_i(clk_edn_i),
        .rst_edn_ni(rst_edn_ni),
        .edn_rnd_o(edn_rnd_o),
        .edn_rnd_i(edn_rnd_i),
        
        .edn_urnd_o(edn_urnd_o),
        .edn_urnd_i(edn_urnd_i)
    );
    
    // Clock Generation
    initial begin 
        clk_i = 0;

        forever begin
            #1 clk_i = ~clk_i;

        end
    end
    
    initial begin 

        cc = 0;
        forever begin
            @(posedge clk_i) ;
            cc = cc + 1;
        end
    end    
    
    initial begin 
        clk_edn_i = 0;
        forever begin
            #1 clk_edn_i = ~clk_edn_i;
        end
    end



    
    // EDN Response Generation
    
    always_ff @ (posedge clk_edn_i)
        begin
            edn_urnd_i = edn_pkg::EDN_RSP_DEFAULT;
            edn_rnd_i = edn_pkg::EDN_RSP_DEFAULT; 
            
            if (edn_urnd_o.edn_req == 1'b1)
                begin
                    edn_urnd_i.edn_ack = edn_urnd_o.edn_req;
                    edn_urnd_i.edn_bus = $urandom();
                end
                
            if (edn_rnd_o.edn_req == 1'b1)
                begin
                    edn_rnd_i.edn_ack = edn_rnd_o.edn_req;
                    edn_rnd_i.edn_bus = $urandom();
                end
             
        end
    
    
    // Tester
    
    initial begin 
        //Inital Bus Signals
        tl_i_d.a_address = 32'h0;
        tl_i_d.a_data = 32'h0;
        tl_i_d.a_mask = 4'hF;
        tl_i_d.a_opcode = tlul_pkg::PutFullData;
        tl_i_d.a_size = 2'b10;
        tl_i_d.a_source = 7'h0;
        tl_i_d.a_valid = 1'b0;
        tl_i_d.a_user = tlul_pkg::TL_A_USER_DEFAULT;
        
        rst_ni = 1;   
        rst_edn_ni = 1;
        #5
        rst_ni = 0;
        rst_edn_ni = 0;
        #5
        rst_ni = 1;   
        rst_edn_ni = 1;
        
        f = $fopen({log_path, "tl_output.txt"},"w");
        
        error_count = 0;
        
        // Header 
        $fwrite(f,"----------------------------------------------------------------\n");
        $fwrite(f,"-- OTBN - RTL - Testbench                                       \n");
        $fwrite(f,"----------------------------------------------------------------\n");
        
        teststate = "Read Registers";
        
        // Read Registers
        for (int i=0 ; i<6 ; i++) begin
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end
        
        // Interrupt Test Register
        read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        teststate = "Run Application";
        // Write Programm to IMEM  
        for (int i=0 ; i<128 ; i++) begin 
            // NOP Instruction
            write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'b10011), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );   
        end
        // ECALL Instruction
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'b1110011), .address(OTBN_IMEM_OFFSET+4*128), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //NOP
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end        
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- MUL256\n");
        $fwrite(f,"----------------------------------------------------------------\n");     
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_mul256.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_mul256.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
        
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        //mul256_expected_result = 
        
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+512), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'h40529766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'hed40926c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'h0622d5ee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'h59b7199e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'h85ab75a5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'h565eff32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'h536bfd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'hdad4a618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'hfa6dc7f2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'h3f2b811b) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10  :   assert (rdbk == 32'h37b795eb) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11  :   assert (rdbk == 32'hea93fcc8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12  :   assert (rdbk == 32'h4cfd63b4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13  :   assert (rdbk == 32'ha0a622d0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14  :   assert (rdbk == 32'h1e3ddfee) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15  :   assert (rdbk == 32'h1066a869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end

        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-PQSR\n");
        $fwrite(f,"----------------------------------------------------------------\n");     
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pqsr.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pqsr.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
        
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        //mul256_expected_result = 
        
        // Read DMEM  
        for (int i=0 ; i<20 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10  :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11  :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12  :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13  :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14  :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15  :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16  :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17  :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18  :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19  :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end
        
        
        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-ADD-SUB\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq-add-sub.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq-add-sub.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
        
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
                
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+512), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'h0000000c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'h0000016a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'h0000000a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'h00000170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'h00000008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'h00000ca4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'h00000006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'h00000cae) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'h00000cfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'h0000083a) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10  :   assert (rdbk == 32'h00000cfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11  :   assert (rdbk == 32'h0000065e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12  :   assert (rdbk == 32'h00000cfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13  :   assert (rdbk == 32'h000003a7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14  :   assert (rdbk == 32'h00000cfd) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15  :   assert (rdbk == 32'h00000051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-MUL\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq-montmul.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq-montmul.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
                
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+512), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'h00000040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'h0000055c) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'h00000031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'h000007da) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'h00000024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'h000004b5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'h00000019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'h00000042) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'h00000bc3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'h000008c1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10  :   assert (rdbk == 32'h000000f5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11  :   assert (rdbk == 32'h00000b67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12  :   assert (rdbk == 32'h00000038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13  :   assert (rdbk == 32'h000003b3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14  :   assert (rdbk == 32'h0000001e) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15  :   assert (rdbk == 32'h00000898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end        


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-BF\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_pq_bf.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_pq_bf.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
                
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+512), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd8023823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd4949942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd5503697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd7227518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4077164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd903461)  else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd2287113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd3389395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd2840445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd1776347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10  :   assert (rdbk == 32'd712249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11  :   assert (rdbk == 32'd8028568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12  :   assert (rdbk == 32'd6964470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13  :   assert (rdbk == 32'd5900372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14  :   assert (rdbk == 32'd4836274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15  :   assert (rdbk == 32'd3772176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
       end     


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-OPT (Dilithium)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_opt_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_opt_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_dilithium = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd8023823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd4949942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd5503697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd7227518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4077164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd903461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd2287113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd3389395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd1447936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd3912035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd3833152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd5335025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd7966085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd8118989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd7144945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd7460296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd8200405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd5651255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd5840697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd2041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd8329041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd2296483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd7624292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd7760084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd6558166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd2463083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd592160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd7596205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd490458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd4570418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd535121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd5905710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd2269315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd25712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd65279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd6056088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd437727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd5437873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd45209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd3628670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd5932184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd4892020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd4400120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd3282855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd5579212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd2040171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd8129297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd3975887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd886499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd5275349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd1715375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd2422113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd503654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2500352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd3475364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd2130347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd7671751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd7706886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd6190567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd1877207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd1880030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd7339689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd5192027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd7408649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd4046506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd6555025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd861568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd5241798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd3351905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd7967553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd8240568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd2908955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd1077579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd7068530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd1063576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd2082141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd1227026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd4901674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd6147942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd4516462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd7784774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd4909015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd2489952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd8055865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd1807242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd3141274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd4210121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd2460839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd6404829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd6055556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd699854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd8144470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd167925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd2815245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd5308330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd7801015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd7301606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd2832490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd6224608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd4233662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd3984450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd6969568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd7183502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd6133025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd3069985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd7499554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd5559452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd7309678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd5405335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd5069329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd3320196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd2451430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd3043243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd3070455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd3966814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd6244424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd2083871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd2186058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd7917105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd5731770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd8357109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd4801012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd3444419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd6442745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd3142318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd4483091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd4065258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd1986703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd8368027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd4615661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd144560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd4178015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd2729052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd7118387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd1224642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd2979664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd2679432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd2620296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd3256914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd7425771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd4495896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd6348741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd6906650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd4571569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd5432259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd4416612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd3304060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd5577029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd3173849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd6062776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd8209741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd1186292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd3076903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd7840971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd2874775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd2013616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd4888110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd5543365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd6149437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd7037817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd2703904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd148603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1178408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd5493962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd2871386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd2394607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd4524768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd626150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd8137948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd2020685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd2930707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd6943539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd3297580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd3309315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd7957803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd3489579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd1101657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd2199934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd2667995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd311407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd4615923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd268380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd7867980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd1165026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd6246419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd7938242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd3436132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd5102358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd1264622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd6021013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd3303556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd104046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd252176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd6426141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd3998553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd918827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd4282041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd2746755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd1284601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd5651462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd6998811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd1817618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd528380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd2525913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd5078866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd8002802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd2110331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd2052914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd155305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd3718478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd5776192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd6905096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd5498888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd7254918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd6047002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd6361152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd915442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd87228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd1281704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd3647397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd8363923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd3451609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd6209053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd1776623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd1128875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd6914893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd4152979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd1018431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd6308070) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd982921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd3563602) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd1283529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd1618324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd1186221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd13008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd759546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd6421303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd5292714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd2462024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd7387771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd7276117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd1343415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd1301221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd977961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd3904031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd193986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd5172786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd1429550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd2425536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd68499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd3777265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd7056830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd6555455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd981963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd8074937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd3279003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-INVNTT-OPT (Dilithium)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_opt_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_opt_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_dilithium_inv = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-OPT (Kyber)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_opt_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_opt_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_kyber = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd2429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd2845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd1865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd1356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd2483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd2197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd2725) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd2668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd2707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd1488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd2194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd1971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd2319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd1075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd3143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd1380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd2718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd1155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd1586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd2874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd1442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd2619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd2169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd2159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd1479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd2634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd2864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd2014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd3200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd1923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd1603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd1732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd1999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd2024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd1094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd2276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd2159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd2187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd1973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd2637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd2158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd2373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd2986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd1482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd1157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd1290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd1057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd2220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd1124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd1019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd2206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd2233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd1376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd2880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd2664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd1960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd1974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd2934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd2679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd2860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd2217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd2897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd3234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd1905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd2306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd2145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd3000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd1378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd2392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd2835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd1685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd1091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd1054) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd2150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd543) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd3192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd2518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd3246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd2277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd2522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd1990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd2637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd3232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd1075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd940) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd2617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd2776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd2606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd2208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd868) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd1949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd2149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd3066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd1896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd2996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd2306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd2463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd1313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd1951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd2999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd1806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd2830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd2104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd1771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd2453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd2605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd1467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd2426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd1985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd2363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd1015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd3120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd3100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd1274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd1919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd1890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd2147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd1961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd1949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd1738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd2772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd1270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd2089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd1051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd2576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd1628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd1735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd3195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd2034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd3195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd2007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd1419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd2334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd2344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd2825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd2523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd2642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd1604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd3280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd1317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd1165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd1532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd3059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd1752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd2052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd1006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd1858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd2336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd1183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd1656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd1668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd2037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd2946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd2184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd1048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd2825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd1363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd1989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd1995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd1551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd2022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd3212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd1591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd1637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd2330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd1625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd2795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd3194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd2717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd3005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd2883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd2594) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd3105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd2502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd2134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd2717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd2303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-INV-OPT (Kyber)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_opt_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_opt_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_kyber_inv = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end

        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-Indirect (Dilithium)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_ind_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_ind_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_dilithium_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd8023823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd4949942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd5503697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd7227518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4077164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd903461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd2287113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd3389395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd1447936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd3912035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd3833152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd5335025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd7966085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd8118989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd7144945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd7460296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd8200405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd5651255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd5840697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd2041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd8329041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd2296483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd7624292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd7760084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd6558166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd2463083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd592160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd7596205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd490458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd4570418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd535121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd5905710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd2269315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd25712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd65279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd6056088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd437727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd5437873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd45209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd3628670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd5932184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd4892020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd4400120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd3282855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd5579212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd2040171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd8129297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd3975887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd886499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd5275349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd1715375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd2422113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd503654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2500352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd3475364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd2130347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd7671751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd7706886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd6190567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd1877207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd1880030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd7339689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd5192027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd7408649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd4046506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd6555025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd861568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd5241798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd3351905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd7967553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd8240568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd2908955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd1077579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd7068530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd1063576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd2082141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd1227026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd4901674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd6147942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd4516462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd7784774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd4909015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd2489952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd8055865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd1807242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd3141274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd4210121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd2460839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd6404829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd6055556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd699854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd8144470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd167925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd2815245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd5308330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd7801015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd7301606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd2832490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd6224608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd4233662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd3984450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd6969568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd7183502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd6133025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd3069985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd7499554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd5559452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd7309678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd5405335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd5069329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd3320196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd2451430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd3043243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd3070455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd3966814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd6244424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd2083871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd2186058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd7917105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd5731770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd8357109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd4801012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd3444419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd6442745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd3142318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd4483091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd4065258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd1986703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd8368027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd4615661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd144560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd4178015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd2729052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd7118387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd1224642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd2979664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd2679432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd2620296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd3256914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd7425771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd4495896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd6348741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd6906650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd4571569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd5432259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd4416612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd3304060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd5577029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd3173849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd6062776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd8209741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd1186292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd3076903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd7840971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd2874775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd2013616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd4888110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd5543365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd6149437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd7037817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd2703904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd148603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1178408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd5493962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd2871386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd2394607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd4524768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd626150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd8137948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd2020685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd2930707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd6943539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd3297580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd3309315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd7957803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd3489579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd1101657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd2199934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd2667995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd311407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd4615923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd268380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd7867980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd1165026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd6246419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd7938242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd3436132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd5102358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd1264622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd6021013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd3303556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd104046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd252176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd6426141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd3998553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd918827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd4282041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd2746755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd1284601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd5651462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd6998811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd1817618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd528380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd2525913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd5078866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd8002802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd2110331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd2052914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd155305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd3718478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd5776192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd6905096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd5498888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd7254918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd6047002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd6361152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd915442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd87228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd1281704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd3647397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd8363923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd3451609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd6209053) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd1776623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd1128875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd6914893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd4152979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd1018431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd6308070) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd982921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd3563602) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd1283529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd1618324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd1186221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd13008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd759546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd6421303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd5292714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd2462024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd7387771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd7276117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd1343415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd1301221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd977961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd3904031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd193986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd5172786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd1429550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd2425536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd68499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd3777265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd7056830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd6555455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd981963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd8074937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd3279003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end

        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-INVNTT Indirect (Dilithium)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_ind_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_ind_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_dilithium_inv_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-Indirect (Kyber)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_ind_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_ind_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_kyber_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd2429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd2845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd1865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd1356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd2483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd2197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd2725) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd2668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd2707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd1488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd2194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd1971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd2319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd1075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd3143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd1380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd2718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd1155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd1586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd2874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd1442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd2619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd2169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd2159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd1479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd2634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd2864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd2014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd3200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd1923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd1603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd1732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd1999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd2024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd1094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd2276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd2159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd2187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd1973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd2637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd2158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd2373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd2986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd1482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd1157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd1290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd1057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd2220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd1124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd1019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd2206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd2233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd1376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd2880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd2664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd1960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd1974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd2934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd2679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd2860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd2217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd2897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd3234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd1905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd2306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd2145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd3000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd1378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd2392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd2835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd1685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd1091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd1054) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd2150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd543) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd3192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd2518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd3246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd2277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd2522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd1990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd2637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd3232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd1075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd940) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd2617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd2776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd2606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd2208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd868) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd1949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd2149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd3066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd1896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd2996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd2306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd2463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd1313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd1951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd2999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd1806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd2830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd2104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd1771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd2453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd2605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd1467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd2426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd1985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd2363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd1015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd3120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd3100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd1274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd1919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd1890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd2147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd1961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd1949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd1738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd2772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd1270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd2089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd1051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd2576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd1628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd1735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd3195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd2034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd3195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd2007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd1419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd2334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd2344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd2825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd2523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd2642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd1604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd3280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd1317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd1165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd1532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd3059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd1752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd2052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd1006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd1858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd2336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd1183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd1656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd1668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd2037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd2946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd2184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd1048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd2825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd1363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd1989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd1995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd1551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd2022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd3212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd1591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd1637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd2330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd1625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd2795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd3194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd2717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd3005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd2883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd2594) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd3105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd2502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd2134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd2717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd2303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-INVNTT Indirect (Kyber)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_ind_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_ind_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_kyber_inv_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+544), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end



        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-Indirect (Falcon-512)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_ind_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_ind_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon512_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<512 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd3478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd8305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd9294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd9394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd6662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd3132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd5560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd3644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd8479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd10395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd9828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd11980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd6723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd6206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd8244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd9116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd8799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd1938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd6517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd3491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd8590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd4573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd3003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd8920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd6129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd1131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd3898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd4583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd1222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd8324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd12266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd4260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd3294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd6324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd6173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd1261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd11311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd5436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd10597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd4052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd6793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd8528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd10528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd9185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd7661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd7160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd11694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd10504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd8452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd5370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd4710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd12110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd4970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd10967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd6398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd5014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd5208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd5550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd4549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd3126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd10965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd7128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd7412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd4171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd6892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd8806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd12189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd10672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd8860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd11349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd10792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd2003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd7810) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd11972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd8697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd11170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd4625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd9323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd2483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd4636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd2111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd8997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd3674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd6965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd2760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd11138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd4506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd2302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd9304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd3880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd5867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd3166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd6674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd6735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd5522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd5118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd8941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd7341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd11250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd10319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd4613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd8373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd11294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd8083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd7760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd5583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd4772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd9982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd1698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd6634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd12261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd8451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd1812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd3451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd4584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd8591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd1331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd1083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd5759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd1373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd7998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd2942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd10805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd5448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd10679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd1256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd7046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd6316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd5909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd9654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd11764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd7025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd7611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd2889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd3751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd6172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd6391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd10611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd7941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd7563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd11079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd4588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd10690) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd3865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd3033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd6576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd4322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd2099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd2549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd4041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd1904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd10519) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd7012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd10196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd7732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd9827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd10792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd4816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd9771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd7304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd8031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd5521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd9032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd1620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd4101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd4303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd5499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd7620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd10736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd8642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd3430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd8118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd8166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd4877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd5304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd7964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd5063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd4584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd9487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd8348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd1734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd2939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd6958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd10013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd3391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd2562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd5609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd4459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd1997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd9743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd5443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd10604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd8722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd8368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd6139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd1825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd5461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd2520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd8926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd11417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd9476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd5541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd11866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd10839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd5724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd1746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd3344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd7852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd8762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd4351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd4068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd11749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd5791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd8103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd7939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd7956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd12126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd6319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd1253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd7230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd8230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd4957) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd5750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd3127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd5092) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd2272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd6433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd6886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd2221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd1973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd8419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd3058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd10731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd8073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd11453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd6766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd6306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd10507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd9219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd4911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd9126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd9699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd3267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd10701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd7238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd4245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd11832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd4718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd4207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd11117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd2188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd1664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd3331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd9465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd6620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd3116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd5582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd9987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd9217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd10393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd7383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd11335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd7057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd2100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd10387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd11657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd3197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd6384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd2256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd7195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd8966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd6343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd9782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd10562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd9990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd6143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd6579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd10741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd8973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd1239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd6050) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd9572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd6346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd10825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd6755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd3082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd6983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd4599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd12059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd1596) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd11382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd2269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd7426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd1130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd6312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd3563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd1410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd10019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd12179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd3443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd11670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd12005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd1256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd1812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd4928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd6449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd10435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd6703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd5618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd7229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd8046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd3908) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd3485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd9999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd8409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd5716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd9779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd10612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd10113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd7087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd2728) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd9673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd10156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd7131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd3222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd5209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd7660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd11592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd4965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd9341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd526) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd8664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd9546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd1536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd3669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd11279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd10845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd11474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd10742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd1391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd6888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd7095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd8088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd8931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd4210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd7058) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd3337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd8259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd10161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd6403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd4704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd4295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd1130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd3146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd12118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd7457) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd12247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd11727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd7340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd5760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd3991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd5890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd3864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd8942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd10354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd8794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd10467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd1009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd2762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd7702) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd4856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd1494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd2156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd4415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd6174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd7215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd10760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd10931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd7300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd3504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd4992) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd10211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd12172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd7585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd4452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd4010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd11778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd2935) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd2829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd1164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd5213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd4509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd10678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd7847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd7948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd5350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd1710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd3253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd3120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd1995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd9425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd7414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd10501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd6805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd7214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd8275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd1856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd5480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd1282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd9736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd2185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd2315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd2226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd11611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd9221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd10590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd7730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd5299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd2380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd5278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd4668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd3233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd1815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd10840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd3421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd5631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd11939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd10708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd4709) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd5447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd3229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd8382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd3826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd7791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd3597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd8338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd10040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd1617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd1191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd3678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd7752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd4197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd3100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd8216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd7443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd6488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd11347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd8865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd1219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd8020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd9646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd9554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd9786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd4045) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end



        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-INVNTT-Indirect (Falcon-512)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_ind_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_ind_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon512_inv_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<512 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd291) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd326) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd328) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd332) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd359) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd367) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd389) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd402) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd434) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd454) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd457) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd460) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd471) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd472) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd475) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd486) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd493) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd505) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd508) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end

        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-NTT-Indirect (Falcon-1024)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_ind_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_ind_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon1024_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<1024 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd5660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd6117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd7575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd11873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd9428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd5469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd5449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd4522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd1799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd9101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd2447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd2339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd9415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd10497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd8616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd11953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd6800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd4677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd1986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd4074) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd2218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd12162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd4464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd1532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd2854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd1578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd8964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd5257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd5925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd5989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd7571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd10995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd2118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd7621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd7308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd5468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd3681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd3495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd4090) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd4201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd1912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd11696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd8473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd6720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd5259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd4886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd10765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd9283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd8861) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd5835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd3145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd9065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd4485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd7885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd1456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd7369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd5525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd2164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd8590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd5722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd3800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd7335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd2802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd6125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd2837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd4174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd4685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd10259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd3785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd8037) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd4567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd4412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd1919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd4691) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd7804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd12106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd1247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd2156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd12180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd8684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd5624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd3071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd5362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd4263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd11224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd10223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd11022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd3029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd9641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd9815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd4010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd8969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd7796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd8428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd11729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd2789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd3569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd9429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd11112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd10591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd6909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd11534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd8143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd6879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd11849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd3624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd11977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd5572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd4337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd10647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd4676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd8126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd5777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd3496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd6375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd1599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd2625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd6154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd2253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd11330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd1184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd1563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd11379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd8515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd8066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd9978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd9988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd10979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd5467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd1401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd6246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd12144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd11241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd3840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd3627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd2936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd7804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd10522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd2546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd8222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd10937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd6775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd12003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd9381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd6279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd4028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd8884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd11513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd3383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd3204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd4385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd1425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd6394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd8439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd5251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd11056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd5140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd4397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd6355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd8557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd12271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd12081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd5791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd2115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd10144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd9144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd5406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd6557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd1557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd2169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd5148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd11654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd6500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd7105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd3905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd11692) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd1038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd5949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd10896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd9340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd1946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd8715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd11530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd8030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd2904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd8968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd5281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd2884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd9286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd6884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd1179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd4934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd3832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd11104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd4933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd6958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd8752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd9820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd9763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd6140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd11737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd8942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd1793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd6901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd6989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd11926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd6004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd1571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd7780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd9774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd3001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd3558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd4020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd7384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd6341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd11712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd9904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd4976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd6409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd10437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd11494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd2325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd1314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd2516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd6846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd8870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd11616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd10635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd5621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd9665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd3189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd9494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd12124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd3016) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd7819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd11466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd11349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd1739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd11141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd8021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd7381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd3759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd11968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd9622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd10046) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd9282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd10881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd1533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd8763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd8758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd2219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd11566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd9225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd10687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd9761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd8476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd8964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd3707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd4916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd1344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd10994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd12098) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd9963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd1833) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd2509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd7758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd1720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd2362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd4802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd9733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd3989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd8666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd9946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd1489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd3299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd5017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd3117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd3431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd5550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd1755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd9313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd1581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd8624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd2355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd9783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd10114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd5276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd10628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd3420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd4101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd10850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd5560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd2035) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd9111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd1100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd4239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd7282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd2398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd2881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd10485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd3639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd11057) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd10188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd1531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd9694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd11605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd2151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd9062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd8570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd9294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd1307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd2452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd11202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd2618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd1703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd7979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd6564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd5309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd4351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd5578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd11815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd4805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd11952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd6307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd11363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd8394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd11307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd5817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd2972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd10746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd3724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd11492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd10863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd5598) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd3117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd5874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd7251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd3264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd6646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd1669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd10024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd11174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd8099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd6001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd8416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd6640) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd10945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd6446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd10580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd4182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd8414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd3368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd10066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd8153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd6099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd1288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd4330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd4394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd1483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd8290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd8113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd12022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd10529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd5638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd7321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd2972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd3571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd3039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd6356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd11008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd6124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd6452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd6926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd8061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd9565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd9356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd3929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd3318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd7265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd4468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd9710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd4803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd4770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd6579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd5071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd2982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd1497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd10113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd4482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd9682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd11039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd7354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd8436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd5665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd2869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd7998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd5718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd9467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd3749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd4956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd8447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd10496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd11803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd10627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd10102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd7682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd1277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd4255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd11229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd7627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd6936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd3027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd2515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd2339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd7313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd2851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd5346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd1481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd8854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd7341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd10075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd3191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd4110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd7843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd10343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd4885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd3771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd11524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd8472) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd2623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd10040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd7927) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd7400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd1585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd11891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd9882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd4854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd3823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd4109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd3192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd5359) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd8327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd4241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd1990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd7253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd2010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd2346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                512   :   assert (rdbk == 32'd4566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                513   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                514   :   assert (rdbk == 32'd997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                515   :   assert (rdbk == 32'd7425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                516   :   assert (rdbk == 32'd2619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                517   :   assert (rdbk == 32'd7567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                518   :   assert (rdbk == 32'd7740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                519   :   assert (rdbk == 32'd1981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                520   :   assert (rdbk == 32'd2357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                521   :   assert (rdbk == 32'd7122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                522   :   assert (rdbk == 32'd9314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                523   :   assert (rdbk == 32'd7314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                524   :   assert (rdbk == 32'd9945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                525   :   assert (rdbk == 32'd4561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                526   :   assert (rdbk == 32'd6611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                527   :   assert (rdbk == 32'd5827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                528   :   assert (rdbk == 32'd4027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                529   :   assert (rdbk == 32'd10647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                530   :   assert (rdbk == 32'd5377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                531   :   assert (rdbk == 32'd4841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                532   :   assert (rdbk == 32'd12169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                533   :   assert (rdbk == 32'd9494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                534   :   assert (rdbk == 32'd8503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                535   :   assert (rdbk == 32'd3571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                536   :   assert (rdbk == 32'd3579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                537   :   assert (rdbk == 32'd1794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                538   :   assert (rdbk == 32'd5911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                539   :   assert (rdbk == 32'd3317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                540   :   assert (rdbk == 32'd1971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                541   :   assert (rdbk == 32'd5904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                542   :   assert (rdbk == 32'd6239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                543   :   assert (rdbk == 32'd2867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                544   :   assert (rdbk == 32'd5239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                545   :   assert (rdbk == 32'd4982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                546   :   assert (rdbk == 32'd267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                547   :   assert (rdbk == 32'd5836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                548   :   assert (rdbk == 32'd10102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                549   :   assert (rdbk == 32'd7324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                550   :   assert (rdbk == 32'd7778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                551   :   assert (rdbk == 32'd3086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                552   :   assert (rdbk == 32'd6484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                553   :   assert (rdbk == 32'd6379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                554   :   assert (rdbk == 32'd4448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                555   :   assert (rdbk == 32'd3228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                556   :   assert (rdbk == 32'd9764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                557   :   assert (rdbk == 32'd7514) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                558   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                559   :   assert (rdbk == 32'd8067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                560   :   assert (rdbk == 32'd7876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                561   :   assert (rdbk == 32'd4961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                562   :   assert (rdbk == 32'd1621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                563   :   assert (rdbk == 32'd1743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                564   :   assert (rdbk == 32'd1743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                565   :   assert (rdbk == 32'd11298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                566   :   assert (rdbk == 32'd2953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                567   :   assert (rdbk == 32'd2871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                568   :   assert (rdbk == 32'd677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                569   :   assert (rdbk == 32'd11476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                570   :   assert (rdbk == 32'd6086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                571   :   assert (rdbk == 32'd8758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                572   :   assert (rdbk == 32'd7723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                573   :   assert (rdbk == 32'd1461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                574   :   assert (rdbk == 32'd6739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                575   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                576   :   assert (rdbk == 32'd9763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                577   :   assert (rdbk == 32'd8570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                578   :   assert (rdbk == 32'd373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                579   :   assert (rdbk == 32'd5812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                580   :   assert (rdbk == 32'd5462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                581   :   assert (rdbk == 32'd746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                582   :   assert (rdbk == 32'd6093) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                583   :   assert (rdbk == 32'd1665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                584   :   assert (rdbk == 32'd5289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                585   :   assert (rdbk == 32'd3846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                586   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                587   :   assert (rdbk == 32'd5182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                588   :   assert (rdbk == 32'd3897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                589   :   assert (rdbk == 32'd7075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                590   :   assert (rdbk == 32'd8970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                591   :   assert (rdbk == 32'd10147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                592   :   assert (rdbk == 32'd5481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                593   :   assert (rdbk == 32'd7667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                594   :   assert (rdbk == 32'd11083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                595   :   assert (rdbk == 32'd3966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                596   :   assert (rdbk == 32'd5283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                597   :   assert (rdbk == 32'd6106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                598   :   assert (rdbk == 32'd4232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                599   :   assert (rdbk == 32'd3084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                600   :   assert (rdbk == 32'd4998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                601   :   assert (rdbk == 32'd1314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                602   :   assert (rdbk == 32'd3636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                603   :   assert (rdbk == 32'd11856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                604   :   assert (rdbk == 32'd8397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                605   :   assert (rdbk == 32'd7463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                606   :   assert (rdbk == 32'd4532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                607   :   assert (rdbk == 32'd5219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                608   :   assert (rdbk == 32'd6511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                609   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                610   :   assert (rdbk == 32'd7849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                611   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                612   :   assert (rdbk == 32'd8807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                613   :   assert (rdbk == 32'd1984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                614   :   assert (rdbk == 32'd8233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                615   :   assert (rdbk == 32'd3761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                616   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                617   :   assert (rdbk == 32'd8529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                618   :   assert (rdbk == 32'd1259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                619   :   assert (rdbk == 32'd9393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                620   :   assert (rdbk == 32'd6759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                621   :   assert (rdbk == 32'd1568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                622   :   assert (rdbk == 32'd5187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                623   :   assert (rdbk == 32'd10634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                624   :   assert (rdbk == 32'd9245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                625   :   assert (rdbk == 32'd3215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                626   :   assert (rdbk == 32'd11521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                627   :   assert (rdbk == 32'd9348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                628   :   assert (rdbk == 32'd8820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                629   :   assert (rdbk == 32'd7716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                630   :   assert (rdbk == 32'd8371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                631   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                632   :   assert (rdbk == 32'd1914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                633   :   assert (rdbk == 32'd2644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                634   :   assert (rdbk == 32'd4243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                635   :   assert (rdbk == 32'd1638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                636   :   assert (rdbk == 32'd2354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                637   :   assert (rdbk == 32'd8712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                638   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                639   :   assert (rdbk == 32'd8305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                640   :   assert (rdbk == 32'd3089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                641   :   assert (rdbk == 32'd8828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                642   :   assert (rdbk == 32'd5856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                643   :   assert (rdbk == 32'd858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                644   :   assert (rdbk == 32'd4477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                645   :   assert (rdbk == 32'd2567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                646   :   assert (rdbk == 32'd10680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                647   :   assert (rdbk == 32'd2467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                648   :   assert (rdbk == 32'd9065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                649   :   assert (rdbk == 32'd7906) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                650   :   assert (rdbk == 32'd2342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                651   :   assert (rdbk == 32'd7567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                652   :   assert (rdbk == 32'd483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                653   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                654   :   assert (rdbk == 32'd257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                655   :   assert (rdbk == 32'd11499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                656   :   assert (rdbk == 32'd6616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                657   :   assert (rdbk == 32'd2870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                658   :   assert (rdbk == 32'd12113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                659   :   assert (rdbk == 32'd5554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                660   :   assert (rdbk == 32'd9996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                661   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                662   :   assert (rdbk == 32'd4630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                663   :   assert (rdbk == 32'd7392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                664   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                665   :   assert (rdbk == 32'd10276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                666   :   assert (rdbk == 32'd11658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                667   :   assert (rdbk == 32'd9667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                668   :   assert (rdbk == 32'd5247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                669   :   assert (rdbk == 32'd10030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                670   :   assert (rdbk == 32'd4814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                671   :   assert (rdbk == 32'd12234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                672   :   assert (rdbk == 32'd6678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                673   :   assert (rdbk == 32'd696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                674   :   assert (rdbk == 32'd10155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                675   :   assert (rdbk == 32'd2740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                676   :   assert (rdbk == 32'd2582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                677   :   assert (rdbk == 32'd11793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                678   :   assert (rdbk == 32'd3161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                679   :   assert (rdbk == 32'd3413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                680   :   assert (rdbk == 32'd10981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                681   :   assert (rdbk == 32'd6885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                682   :   assert (rdbk == 32'd11440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                683   :   assert (rdbk == 32'd511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                684   :   assert (rdbk == 32'd3726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                685   :   assert (rdbk == 32'd3649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                686   :   assert (rdbk == 32'd11686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                687   :   assert (rdbk == 32'd10147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                688   :   assert (rdbk == 32'd5641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                689   :   assert (rdbk == 32'd12152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                690   :   assert (rdbk == 32'd10550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                691   :   assert (rdbk == 32'd11544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                692   :   assert (rdbk == 32'd8848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                693   :   assert (rdbk == 32'd381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                694   :   assert (rdbk == 32'd979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                695   :   assert (rdbk == 32'd5847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                696   :   assert (rdbk == 32'd11590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                697   :   assert (rdbk == 32'd7655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                698   :   assert (rdbk == 32'd951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                699   :   assert (rdbk == 32'd8417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                700   :   assert (rdbk == 32'd9096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                701   :   assert (rdbk == 32'd10900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                702   :   assert (rdbk == 32'd8126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                703   :   assert (rdbk == 32'd2962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                704   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                705   :   assert (rdbk == 32'd10767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                706   :   assert (rdbk == 32'd8559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                707   :   assert (rdbk == 32'd9181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                708   :   assert (rdbk == 32'd12232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                709   :   assert (rdbk == 32'd11077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                710   :   assert (rdbk == 32'd4563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                711   :   assert (rdbk == 32'd12232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                712   :   assert (rdbk == 32'd275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                713   :   assert (rdbk == 32'd5106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                714   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                715   :   assert (rdbk == 32'd9180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                716   :   assert (rdbk == 32'd1032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                717   :   assert (rdbk == 32'd11960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                718   :   assert (rdbk == 32'd5312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                719   :   assert (rdbk == 32'd419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                720   :   assert (rdbk == 32'd7311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                721   :   assert (rdbk == 32'd10911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                722   :   assert (rdbk == 32'd11165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                723   :   assert (rdbk == 32'd4435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                724   :   assert (rdbk == 32'd3750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                725   :   assert (rdbk == 32'd4521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                726   :   assert (rdbk == 32'd11119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                727   :   assert (rdbk == 32'd4012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                728   :   assert (rdbk == 32'd5070) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                729   :   assert (rdbk == 32'd6650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                730   :   assert (rdbk == 32'd10616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                731   :   assert (rdbk == 32'd2061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                732   :   assert (rdbk == 32'd10680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                733   :   assert (rdbk == 32'd6930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                734   :   assert (rdbk == 32'd7706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                735   :   assert (rdbk == 32'd6985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                736   :   assert (rdbk == 32'd6417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                737   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                738   :   assert (rdbk == 32'd7287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                739   :   assert (rdbk == 32'd10529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                740   :   assert (rdbk == 32'd7219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                741   :   assert (rdbk == 32'd1634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                742   :   assert (rdbk == 32'd5891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                743   :   assert (rdbk == 32'd2208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                744   :   assert (rdbk == 32'd11568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                745   :   assert (rdbk == 32'd6189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                746   :   assert (rdbk == 32'd2119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                747   :   assert (rdbk == 32'd5895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                748   :   assert (rdbk == 32'd7544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                749   :   assert (rdbk == 32'd991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                750   :   assert (rdbk == 32'd4339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                751   :   assert (rdbk == 32'd3685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                752   :   assert (rdbk == 32'd2121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                753   :   assert (rdbk == 32'd8753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                754   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                755   :   assert (rdbk == 32'd6846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                756   :   assert (rdbk == 32'd5681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                757   :   assert (rdbk == 32'd6881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                758   :   assert (rdbk == 32'd9477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                759   :   assert (rdbk == 32'd10942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                760   :   assert (rdbk == 32'd9380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                761   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                762   :   assert (rdbk == 32'd5278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                763   :   assert (rdbk == 32'd3582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                764   :   assert (rdbk == 32'd7958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                765   :   assert (rdbk == 32'd6407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                766   :   assert (rdbk == 32'd9539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                767   :   assert (rdbk == 32'd4727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                768   :   assert (rdbk == 32'd919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                769   :   assert (rdbk == 32'd816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                770   :   assert (rdbk == 32'd10272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                771   :   assert (rdbk == 32'd10916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                772   :   assert (rdbk == 32'd1701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                773   :   assert (rdbk == 32'd4988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                774   :   assert (rdbk == 32'd6354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                775   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                776   :   assert (rdbk == 32'd11504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                777   :   assert (rdbk == 32'd8218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                778   :   assert (rdbk == 32'd11557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                779   :   assert (rdbk == 32'd9012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                780   :   assert (rdbk == 32'd9003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                781   :   assert (rdbk == 32'd10068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                782   :   assert (rdbk == 32'd7205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                783   :   assert (rdbk == 32'd2845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                784   :   assert (rdbk == 32'd8731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                785   :   assert (rdbk == 32'd8122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                786   :   assert (rdbk == 32'd4167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                787   :   assert (rdbk == 32'd6881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                788   :   assert (rdbk == 32'd9430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                789   :   assert (rdbk == 32'd11557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                790   :   assert (rdbk == 32'd9823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                791   :   assert (rdbk == 32'd10649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                792   :   assert (rdbk == 32'd7192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                793   :   assert (rdbk == 32'd2355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                794   :   assert (rdbk == 32'd448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                795   :   assert (rdbk == 32'd3547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                796   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                797   :   assert (rdbk == 32'd5307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                798   :   assert (rdbk == 32'd3361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                799   :   assert (rdbk == 32'd6225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                800   :   assert (rdbk == 32'd11565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                801   :   assert (rdbk == 32'd7951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                802   :   assert (rdbk == 32'd4476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                803   :   assert (rdbk == 32'd10055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                804   :   assert (rdbk == 32'd4380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                805   :   assert (rdbk == 32'd1212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                806   :   assert (rdbk == 32'd9560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                807   :   assert (rdbk == 32'd6651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                808   :   assert (rdbk == 32'd3403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                809   :   assert (rdbk == 32'd5777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                810   :   assert (rdbk == 32'd7708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                811   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                812   :   assert (rdbk == 32'd5364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                813   :   assert (rdbk == 32'd3352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                814   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                815   :   assert (rdbk == 32'd5304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                816   :   assert (rdbk == 32'd10540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                817   :   assert (rdbk == 32'd10257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                818   :   assert (rdbk == 32'd1768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                819   :   assert (rdbk == 32'd7014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                820   :   assert (rdbk == 32'd1921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                821   :   assert (rdbk == 32'd10607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                822   :   assert (rdbk == 32'd9384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                823   :   assert (rdbk == 32'd10657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                824   :   assert (rdbk == 32'd10948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                825   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                826   :   assert (rdbk == 32'd5291) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                827   :   assert (rdbk == 32'd7395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                828   :   assert (rdbk == 32'd5916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                829   :   assert (rdbk == 32'd9887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                830   :   assert (rdbk == 32'd417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                831   :   assert (rdbk == 32'd5760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                832   :   assert (rdbk == 32'd6027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                833   :   assert (rdbk == 32'd1562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                834   :   assert (rdbk == 32'd4114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                835   :   assert (rdbk == 32'd6746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                836   :   assert (rdbk == 32'd9680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                837   :   assert (rdbk == 32'd6129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                838   :   assert (rdbk == 32'd8003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                839   :   assert (rdbk == 32'd5233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                840   :   assert (rdbk == 32'd1495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                841   :   assert (rdbk == 32'd4645) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                842   :   assert (rdbk == 32'd4752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                843   :   assert (rdbk == 32'd11487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                844   :   assert (rdbk == 32'd755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                845   :   assert (rdbk == 32'd8890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                846   :   assert (rdbk == 32'd4126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                847   :   assert (rdbk == 32'd5381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                848   :   assert (rdbk == 32'd4723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                849   :   assert (rdbk == 32'd1837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                850   :   assert (rdbk == 32'd11599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                851   :   assert (rdbk == 32'd5527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                852   :   assert (rdbk == 32'd1137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                853   :   assert (rdbk == 32'd11898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                854   :   assert (rdbk == 32'd3503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                855   :   assert (rdbk == 32'd5542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                856   :   assert (rdbk == 32'd5065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                857   :   assert (rdbk == 32'd2144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                858   :   assert (rdbk == 32'd2351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                859   :   assert (rdbk == 32'd6358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                860   :   assert (rdbk == 32'd11126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                861   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                862   :   assert (rdbk == 32'd2742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                863   :   assert (rdbk == 32'd5199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                864   :   assert (rdbk == 32'd5720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                865   :   assert (rdbk == 32'd9439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                866   :   assert (rdbk == 32'd10943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                867   :   assert (rdbk == 32'd10208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                868   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                869   :   assert (rdbk == 32'd8666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                870   :   assert (rdbk == 32'd11895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                871   :   assert (rdbk == 32'd1073) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                872   :   assert (rdbk == 32'd1795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                873   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                874   :   assert (rdbk == 32'd8664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                875   :   assert (rdbk == 32'd2892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                876   :   assert (rdbk == 32'd6747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                877   :   assert (rdbk == 32'd2029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                878   :   assert (rdbk == 32'd6024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                879   :   assert (rdbk == 32'd11867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                880   :   assert (rdbk == 32'd7355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                881   :   assert (rdbk == 32'd5503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                882   :   assert (rdbk == 32'd1441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                883   :   assert (rdbk == 32'd7953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                884   :   assert (rdbk == 32'd6012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                885   :   assert (rdbk == 32'd2726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                886   :   assert (rdbk == 32'd6583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                887   :   assert (rdbk == 32'd7731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                888   :   assert (rdbk == 32'd3015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                889   :   assert (rdbk == 32'd7420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                890   :   assert (rdbk == 32'd1902) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                891   :   assert (rdbk == 32'd11923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                892   :   assert (rdbk == 32'd10773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                893   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                894   :   assert (rdbk == 32'd11656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                895   :   assert (rdbk == 32'd3257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                896   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                897   :   assert (rdbk == 32'd10357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                898   :   assert (rdbk == 32'd268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                899   :   assert (rdbk == 32'd8695) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                900   :   assert (rdbk == 32'd8445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                901   :   assert (rdbk == 32'd1268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                902   :   assert (rdbk == 32'd11945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                903   :   assert (rdbk == 32'd8144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                904   :   assert (rdbk == 32'd11254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                905   :   assert (rdbk == 32'd10123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                906   :   assert (rdbk == 32'd7628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                907   :   assert (rdbk == 32'd5082) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                908   :   assert (rdbk == 32'd8264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                909   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                910   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                911   :   assert (rdbk == 32'd7201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                912   :   assert (rdbk == 32'd6158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                913   :   assert (rdbk == 32'd1825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                914   :   assert (rdbk == 32'd6382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                915   :   assert (rdbk == 32'd2766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                916   :   assert (rdbk == 32'd9797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                917   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                918   :   assert (rdbk == 32'd7320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                919   :   assert (rdbk == 32'd3460) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                920   :   assert (rdbk == 32'd5849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                921   :   assert (rdbk == 32'd4764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                922   :   assert (rdbk == 32'd4496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                923   :   assert (rdbk == 32'd1590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                924   :   assert (rdbk == 32'd10785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                925   :   assert (rdbk == 32'd7963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                926   :   assert (rdbk == 32'd9156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                927   :   assert (rdbk == 32'd3823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                928   :   assert (rdbk == 32'd8440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                929   :   assert (rdbk == 32'd7431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                930   :   assert (rdbk == 32'd11985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                931   :   assert (rdbk == 32'd1813) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                932   :   assert (rdbk == 32'd8294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                933   :   assert (rdbk == 32'd333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                934   :   assert (rdbk == 32'd2819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                935   :   assert (rdbk == 32'd1315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                936   :   assert (rdbk == 32'd5125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                937   :   assert (rdbk == 32'd10219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                938   :   assert (rdbk == 32'd3029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                939   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                940   :   assert (rdbk == 32'd1107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                941   :   assert (rdbk == 32'd4023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                942   :   assert (rdbk == 32'd10019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                943   :   assert (rdbk == 32'd12223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                944   :   assert (rdbk == 32'd6310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                945   :   assert (rdbk == 32'd12054) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                946   :   assert (rdbk == 32'd7680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                947   :   assert (rdbk == 32'd10999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                948   :   assert (rdbk == 32'd7734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                949   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                950   :   assert (rdbk == 32'd2587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                951   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                952   :   assert (rdbk == 32'd3000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                953   :   assert (rdbk == 32'd4632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                954   :   assert (rdbk == 32'd8608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                955   :   assert (rdbk == 32'd8859) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                956   :   assert (rdbk == 32'd2429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                957   :   assert (rdbk == 32'd11232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                958   :   assert (rdbk == 32'd2622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                959   :   assert (rdbk == 32'd6641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                960   :   assert (rdbk == 32'd4520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                961   :   assert (rdbk == 32'd9522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                962   :   assert (rdbk == 32'd4442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                963   :   assert (rdbk == 32'd7312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                964   :   assert (rdbk == 32'd3089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                965   :   assert (rdbk == 32'd7560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                966   :   assert (rdbk == 32'd10622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                967   :   assert (rdbk == 32'd6280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                968   :   assert (rdbk == 32'd5464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                969   :   assert (rdbk == 32'd4180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                970   :   assert (rdbk == 32'd7974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                971   :   assert (rdbk == 32'd2365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                972   :   assert (rdbk == 32'd2414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                973   :   assert (rdbk == 32'd872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                974   :   assert (rdbk == 32'd656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                975   :   assert (rdbk == 32'd8956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                976   :   assert (rdbk == 32'd6630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                977   :   assert (rdbk == 32'd8287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                978   :   assert (rdbk == 32'd10527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                979   :   assert (rdbk == 32'd11047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                980   :   assert (rdbk == 32'd4752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                981   :   assert (rdbk == 32'd8244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                982   :   assert (rdbk == 32'd9886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                983   :   assert (rdbk == 32'd4409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                984   :   assert (rdbk == 32'd2404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                985   :   assert (rdbk == 32'd12024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                986   :   assert (rdbk == 32'd1892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                987   :   assert (rdbk == 32'd8732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                988   :   assert (rdbk == 32'd2897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                989   :   assert (rdbk == 32'd4841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                990   :   assert (rdbk == 32'd4950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                991   :   assert (rdbk == 32'd12236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                992   :   assert (rdbk == 32'd6976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                993   :   assert (rdbk == 32'd2983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                994   :   assert (rdbk == 32'd2006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                995   :   assert (rdbk == 32'd11065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                996   :   assert (rdbk == 32'd9029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                997   :   assert (rdbk == 32'd4067) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                998   :   assert (rdbk == 32'd3719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                999   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1000   :   assert (rdbk == 32'd5194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1001   :   assert (rdbk == 32'd7619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1002   :   assert (rdbk == 32'd2080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1003   :   assert (rdbk == 32'd8898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1004   :   assert (rdbk == 32'd2821) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1005   :   assert (rdbk == 32'd6363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1006   :   assert (rdbk == 32'd5697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1007   :   assert (rdbk == 32'd3777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1008   :   assert (rdbk == 32'd9416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1009   :   assert (rdbk == 32'd534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1010   :   assert (rdbk == 32'd9793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1011   :   assert (rdbk == 32'd9051) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1012   :   assert (rdbk == 32'd6480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1013   :   assert (rdbk == 32'd7324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1014   :   assert (rdbk == 32'd11620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1015   :   assert (rdbk == 32'd7411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1016   :   assert (rdbk == 32'd11198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1017   :   assert (rdbk == 32'd1298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1018   :   assert (rdbk == 32'd1011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1019   :   assert (rdbk == 32'd10767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1020   :   assert (rdbk == 32'd10026) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1021   :   assert (rdbk == 32'd4756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1022   :   assert (rdbk == 32'd3028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1023   :   assert (rdbk == 32'd4733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end



        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- PQ-INVNTT-Indirect (Falcon-1024)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_ntt_inv_ind_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_ntt_inv_ind_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon1024_inv_indirect = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<1024 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+192), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd2) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd3) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd5) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd6) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd7) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd8) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd10) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd11) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd13) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd14) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd18) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd19) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd20) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd21) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd22) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd23) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd24) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd26) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd27) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd29) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd30) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd31) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd33) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd34) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd35) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd37) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd38) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd39) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd41) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd43) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd44) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd45) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd46) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd47) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd48) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd50) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd52) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd53) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd54) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd55) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd56) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd57) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd58) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd60) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd63) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd65) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd66) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd67) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd68) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd69) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd70) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd72) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd73) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd74) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd75) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd76) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd77) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd78) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd79) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd80) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd82) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd83) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd86) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd87) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd88) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd89) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd90) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd91) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd92) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd93) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd94) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd95) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd97) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd98) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd99) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd103) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd109) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd114) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd131) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd140) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd147) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd148) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd149) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd150) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd151) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd153) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd162) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd172) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd174) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd175) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd178) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd190) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd192) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd194) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd203) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd212) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd213) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd219) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd230) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd246) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd252) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd257) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd258) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd261) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd266) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd275) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd287) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd291) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd293) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd294) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd298) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd299) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd302) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd303) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd305) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd306) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd307) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd308) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd314) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd315) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd317) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd326) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd328) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd332) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd334) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd339) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd340) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd341) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd345) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd347) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd350) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd353) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd359) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd367) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd370) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd387) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd389) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd392) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd399) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd402) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd406) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd407) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd411) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd412) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd419) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd421) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd425) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd432) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd433) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd434) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd437) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd445) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd454) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd457) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd460) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd466) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd468) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd471) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd472) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd475) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd478) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd479) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd486) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd490) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd493) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd497) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd498) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd501) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd505) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd506) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd508) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                512   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                513   :   assert (rdbk == 32'd513) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                514   :   assert (rdbk == 32'd514) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                515   :   assert (rdbk == 32'd515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                516   :   assert (rdbk == 32'd516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                517   :   assert (rdbk == 32'd517) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                518   :   assert (rdbk == 32'd518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                519   :   assert (rdbk == 32'd519) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                520   :   assert (rdbk == 32'd520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                521   :   assert (rdbk == 32'd521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                522   :   assert (rdbk == 32'd522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                523   :   assert (rdbk == 32'd523) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                524   :   assert (rdbk == 32'd524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                525   :   assert (rdbk == 32'd525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                526   :   assert (rdbk == 32'd526) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                527   :   assert (rdbk == 32'd527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                528   :   assert (rdbk == 32'd528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                529   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                530   :   assert (rdbk == 32'd530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                531   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                532   :   assert (rdbk == 32'd532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                533   :   assert (rdbk == 32'd533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                534   :   assert (rdbk == 32'd534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                535   :   assert (rdbk == 32'd535) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                536   :   assert (rdbk == 32'd536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                537   :   assert (rdbk == 32'd537) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                538   :   assert (rdbk == 32'd538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                539   :   assert (rdbk == 32'd539) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                540   :   assert (rdbk == 32'd540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                541   :   assert (rdbk == 32'd541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                542   :   assert (rdbk == 32'd542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                543   :   assert (rdbk == 32'd543) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                544   :   assert (rdbk == 32'd544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                545   :   assert (rdbk == 32'd545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                546   :   assert (rdbk == 32'd546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                547   :   assert (rdbk == 32'd547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                548   :   assert (rdbk == 32'd548) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                549   :   assert (rdbk == 32'd549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                550   :   assert (rdbk == 32'd550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                551   :   assert (rdbk == 32'd551) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                552   :   assert (rdbk == 32'd552) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                553   :   assert (rdbk == 32'd553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                554   :   assert (rdbk == 32'd554) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                555   :   assert (rdbk == 32'd555) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                556   :   assert (rdbk == 32'd556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                557   :   assert (rdbk == 32'd557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                558   :   assert (rdbk == 32'd558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                559   :   assert (rdbk == 32'd559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                560   :   assert (rdbk == 32'd560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                561   :   assert (rdbk == 32'd561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                562   :   assert (rdbk == 32'd562) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                563   :   assert (rdbk == 32'd563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                564   :   assert (rdbk == 32'd564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                565   :   assert (rdbk == 32'd565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                566   :   assert (rdbk == 32'd566) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                567   :   assert (rdbk == 32'd567) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                568   :   assert (rdbk == 32'd568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                569   :   assert (rdbk == 32'd569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                570   :   assert (rdbk == 32'd570) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                571   :   assert (rdbk == 32'd571) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                572   :   assert (rdbk == 32'd572) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                573   :   assert (rdbk == 32'd573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                574   :   assert (rdbk == 32'd574) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                575   :   assert (rdbk == 32'd575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                576   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                577   :   assert (rdbk == 32'd577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                578   :   assert (rdbk == 32'd578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                579   :   assert (rdbk == 32'd579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                580   :   assert (rdbk == 32'd580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                581   :   assert (rdbk == 32'd581) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                582   :   assert (rdbk == 32'd582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                583   :   assert (rdbk == 32'd583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                584   :   assert (rdbk == 32'd584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                585   :   assert (rdbk == 32'd585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                586   :   assert (rdbk == 32'd586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                587   :   assert (rdbk == 32'd587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                588   :   assert (rdbk == 32'd588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                589   :   assert (rdbk == 32'd589) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                590   :   assert (rdbk == 32'd590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                591   :   assert (rdbk == 32'd591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                592   :   assert (rdbk == 32'd592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                593   :   assert (rdbk == 32'd593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                594   :   assert (rdbk == 32'd594) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                595   :   assert (rdbk == 32'd595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                596   :   assert (rdbk == 32'd596) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                597   :   assert (rdbk == 32'd597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                598   :   assert (rdbk == 32'd598) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                599   :   assert (rdbk == 32'd599) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                600   :   assert (rdbk == 32'd600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                601   :   assert (rdbk == 32'd601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                602   :   assert (rdbk == 32'd602) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                603   :   assert (rdbk == 32'd603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                604   :   assert (rdbk == 32'd604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                605   :   assert (rdbk == 32'd605) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                606   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                607   :   assert (rdbk == 32'd607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                608   :   assert (rdbk == 32'd608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                609   :   assert (rdbk == 32'd609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                610   :   assert (rdbk == 32'd610) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                611   :   assert (rdbk == 32'd611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                612   :   assert (rdbk == 32'd612) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                613   :   assert (rdbk == 32'd613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                614   :   assert (rdbk == 32'd614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                615   :   assert (rdbk == 32'd615) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                616   :   assert (rdbk == 32'd616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                617   :   assert (rdbk == 32'd617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                618   :   assert (rdbk == 32'd618) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                619   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                620   :   assert (rdbk == 32'd620) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                621   :   assert (rdbk == 32'd621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                622   :   assert (rdbk == 32'd622) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                623   :   assert (rdbk == 32'd623) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                624   :   assert (rdbk == 32'd624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                625   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                626   :   assert (rdbk == 32'd626) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                627   :   assert (rdbk == 32'd627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                628   :   assert (rdbk == 32'd628) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                629   :   assert (rdbk == 32'd629) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                630   :   assert (rdbk == 32'd630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                631   :   assert (rdbk == 32'd631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                632   :   assert (rdbk == 32'd632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                633   :   assert (rdbk == 32'd633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                634   :   assert (rdbk == 32'd634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                635   :   assert (rdbk == 32'd635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                636   :   assert (rdbk == 32'd636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                637   :   assert (rdbk == 32'd637) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                638   :   assert (rdbk == 32'd638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                639   :   assert (rdbk == 32'd639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                640   :   assert (rdbk == 32'd640) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                641   :   assert (rdbk == 32'd641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                642   :   assert (rdbk == 32'd642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                643   :   assert (rdbk == 32'd643) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                644   :   assert (rdbk == 32'd644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                645   :   assert (rdbk == 32'd645) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                646   :   assert (rdbk == 32'd646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                647   :   assert (rdbk == 32'd647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                648   :   assert (rdbk == 32'd648) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                649   :   assert (rdbk == 32'd649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                650   :   assert (rdbk == 32'd650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                651   :   assert (rdbk == 32'd651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                652   :   assert (rdbk == 32'd652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                653   :   assert (rdbk == 32'd653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                654   :   assert (rdbk == 32'd654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                655   :   assert (rdbk == 32'd655) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                656   :   assert (rdbk == 32'd656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                657   :   assert (rdbk == 32'd657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                658   :   assert (rdbk == 32'd658) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                659   :   assert (rdbk == 32'd659) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                660   :   assert (rdbk == 32'd660) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                661   :   assert (rdbk == 32'd661) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                662   :   assert (rdbk == 32'd662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                663   :   assert (rdbk == 32'd663) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                664   :   assert (rdbk == 32'd664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                665   :   assert (rdbk == 32'd665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                666   :   assert (rdbk == 32'd666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                667   :   assert (rdbk == 32'd667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                668   :   assert (rdbk == 32'd668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                669   :   assert (rdbk == 32'd669) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                670   :   assert (rdbk == 32'd670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                671   :   assert (rdbk == 32'd671) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                672   :   assert (rdbk == 32'd672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                673   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                674   :   assert (rdbk == 32'd674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                675   :   assert (rdbk == 32'd675) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                676   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                677   :   assert (rdbk == 32'd677) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                678   :   assert (rdbk == 32'd678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                679   :   assert (rdbk == 32'd679) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                680   :   assert (rdbk == 32'd680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                681   :   assert (rdbk == 32'd681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                682   :   assert (rdbk == 32'd682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                683   :   assert (rdbk == 32'd683) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                684   :   assert (rdbk == 32'd684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                685   :   assert (rdbk == 32'd685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                686   :   assert (rdbk == 32'd686) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                687   :   assert (rdbk == 32'd687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                688   :   assert (rdbk == 32'd688) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                689   :   assert (rdbk == 32'd689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                690   :   assert (rdbk == 32'd690) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                691   :   assert (rdbk == 32'd691) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                692   :   assert (rdbk == 32'd692) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                693   :   assert (rdbk == 32'd693) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                694   :   assert (rdbk == 32'd694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                695   :   assert (rdbk == 32'd695) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                696   :   assert (rdbk == 32'd696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                697   :   assert (rdbk == 32'd697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                698   :   assert (rdbk == 32'd698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                699   :   assert (rdbk == 32'd699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                700   :   assert (rdbk == 32'd700) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                701   :   assert (rdbk == 32'd701) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                702   :   assert (rdbk == 32'd702) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                703   :   assert (rdbk == 32'd703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                704   :   assert (rdbk == 32'd704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                705   :   assert (rdbk == 32'd705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                706   :   assert (rdbk == 32'd706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                707   :   assert (rdbk == 32'd707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                708   :   assert (rdbk == 32'd708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                709   :   assert (rdbk == 32'd709) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                710   :   assert (rdbk == 32'd710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                711   :   assert (rdbk == 32'd711) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                712   :   assert (rdbk == 32'd712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                713   :   assert (rdbk == 32'd713) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                714   :   assert (rdbk == 32'd714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                715   :   assert (rdbk == 32'd715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                716   :   assert (rdbk == 32'd716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                717   :   assert (rdbk == 32'd717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                718   :   assert (rdbk == 32'd718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                719   :   assert (rdbk == 32'd719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                720   :   assert (rdbk == 32'd720) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                721   :   assert (rdbk == 32'd721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                722   :   assert (rdbk == 32'd722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                723   :   assert (rdbk == 32'd723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                724   :   assert (rdbk == 32'd724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                725   :   assert (rdbk == 32'd725) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                726   :   assert (rdbk == 32'd726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                727   :   assert (rdbk == 32'd727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                728   :   assert (rdbk == 32'd728) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                729   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                730   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                731   :   assert (rdbk == 32'd731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                732   :   assert (rdbk == 32'd732) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                733   :   assert (rdbk == 32'd733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                734   :   assert (rdbk == 32'd734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                735   :   assert (rdbk == 32'd735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                736   :   assert (rdbk == 32'd736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                737   :   assert (rdbk == 32'd737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                738   :   assert (rdbk == 32'd738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                739   :   assert (rdbk == 32'd739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                740   :   assert (rdbk == 32'd740) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                741   :   assert (rdbk == 32'd741) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                742   :   assert (rdbk == 32'd742) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                743   :   assert (rdbk == 32'd743) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                744   :   assert (rdbk == 32'd744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                745   :   assert (rdbk == 32'd745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                746   :   assert (rdbk == 32'd746) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                747   :   assert (rdbk == 32'd747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                748   :   assert (rdbk == 32'd748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                749   :   assert (rdbk == 32'd749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                750   :   assert (rdbk == 32'd750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                751   :   assert (rdbk == 32'd751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                752   :   assert (rdbk == 32'd752) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                753   :   assert (rdbk == 32'd753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                754   :   assert (rdbk == 32'd754) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                755   :   assert (rdbk == 32'd755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                756   :   assert (rdbk == 32'd756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                757   :   assert (rdbk == 32'd757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                758   :   assert (rdbk == 32'd758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                759   :   assert (rdbk == 32'd759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                760   :   assert (rdbk == 32'd760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                761   :   assert (rdbk == 32'd761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                762   :   assert (rdbk == 32'd762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                763   :   assert (rdbk == 32'd763) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                764   :   assert (rdbk == 32'd764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                765   :   assert (rdbk == 32'd765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                766   :   assert (rdbk == 32'd766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                767   :   assert (rdbk == 32'd767) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                768   :   assert (rdbk == 32'd768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                769   :   assert (rdbk == 32'd769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                770   :   assert (rdbk == 32'd770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                771   :   assert (rdbk == 32'd771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                772   :   assert (rdbk == 32'd772) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                773   :   assert (rdbk == 32'd773) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                774   :   assert (rdbk == 32'd774) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                775   :   assert (rdbk == 32'd775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                776   :   assert (rdbk == 32'd776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                777   :   assert (rdbk == 32'd777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                778   :   assert (rdbk == 32'd778) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                779   :   assert (rdbk == 32'd779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                780   :   assert (rdbk == 32'd780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                781   :   assert (rdbk == 32'd781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                782   :   assert (rdbk == 32'd782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                783   :   assert (rdbk == 32'd783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                784   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                785   :   assert (rdbk == 32'd785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                786   :   assert (rdbk == 32'd786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                787   :   assert (rdbk == 32'd787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                788   :   assert (rdbk == 32'd788) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                789   :   assert (rdbk == 32'd789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                790   :   assert (rdbk == 32'd790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                791   :   assert (rdbk == 32'd791) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                792   :   assert (rdbk == 32'd792) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                793   :   assert (rdbk == 32'd793) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                794   :   assert (rdbk == 32'd794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                795   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                796   :   assert (rdbk == 32'd796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                797   :   assert (rdbk == 32'd797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                798   :   assert (rdbk == 32'd798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                799   :   assert (rdbk == 32'd799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                800   :   assert (rdbk == 32'd800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                801   :   assert (rdbk == 32'd801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                802   :   assert (rdbk == 32'd802) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                803   :   assert (rdbk == 32'd803) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                804   :   assert (rdbk == 32'd804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                805   :   assert (rdbk == 32'd805) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                806   :   assert (rdbk == 32'd806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                807   :   assert (rdbk == 32'd807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                808   :   assert (rdbk == 32'd808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                809   :   assert (rdbk == 32'd809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                810   :   assert (rdbk == 32'd810) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                811   :   assert (rdbk == 32'd811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                812   :   assert (rdbk == 32'd812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                813   :   assert (rdbk == 32'd813) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                814   :   assert (rdbk == 32'd814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                815   :   assert (rdbk == 32'd815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                816   :   assert (rdbk == 32'd816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                817   :   assert (rdbk == 32'd817) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                818   :   assert (rdbk == 32'd818) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                819   :   assert (rdbk == 32'd819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                820   :   assert (rdbk == 32'd820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                821   :   assert (rdbk == 32'd821) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                822   :   assert (rdbk == 32'd822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                823   :   assert (rdbk == 32'd823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                824   :   assert (rdbk == 32'd824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                825   :   assert (rdbk == 32'd825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                826   :   assert (rdbk == 32'd826) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                827   :   assert (rdbk == 32'd827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                828   :   assert (rdbk == 32'd828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                829   :   assert (rdbk == 32'd829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                830   :   assert (rdbk == 32'd830) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                831   :   assert (rdbk == 32'd831) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                832   :   assert (rdbk == 32'd832) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                833   :   assert (rdbk == 32'd833) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                834   :   assert (rdbk == 32'd834) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                835   :   assert (rdbk == 32'd835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                836   :   assert (rdbk == 32'd836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                837   :   assert (rdbk == 32'd837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                838   :   assert (rdbk == 32'd838) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                839   :   assert (rdbk == 32'd839) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                840   :   assert (rdbk == 32'd840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                841   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                842   :   assert (rdbk == 32'd842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                843   :   assert (rdbk == 32'd843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                844   :   assert (rdbk == 32'd844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                845   :   assert (rdbk == 32'd845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                846   :   assert (rdbk == 32'd846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                847   :   assert (rdbk == 32'd847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                848   :   assert (rdbk == 32'd848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                849   :   assert (rdbk == 32'd849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                850   :   assert (rdbk == 32'd850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                851   :   assert (rdbk == 32'd851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                852   :   assert (rdbk == 32'd852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                853   :   assert (rdbk == 32'd853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                854   :   assert (rdbk == 32'd854) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                855   :   assert (rdbk == 32'd855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                856   :   assert (rdbk == 32'd856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                857   :   assert (rdbk == 32'd857) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                858   :   assert (rdbk == 32'd858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                859   :   assert (rdbk == 32'd859) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                860   :   assert (rdbk == 32'd860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                861   :   assert (rdbk == 32'd861) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                862   :   assert (rdbk == 32'd862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                863   :   assert (rdbk == 32'd863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                864   :   assert (rdbk == 32'd864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                865   :   assert (rdbk == 32'd865) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                866   :   assert (rdbk == 32'd866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                867   :   assert (rdbk == 32'd867) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                868   :   assert (rdbk == 32'd868) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                869   :   assert (rdbk == 32'd869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                870   :   assert (rdbk == 32'd870) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                871   :   assert (rdbk == 32'd871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                872   :   assert (rdbk == 32'd872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                873   :   assert (rdbk == 32'd873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                874   :   assert (rdbk == 32'd874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                875   :   assert (rdbk == 32'd875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                876   :   assert (rdbk == 32'd876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                877   :   assert (rdbk == 32'd877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                878   :   assert (rdbk == 32'd878) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                879   :   assert (rdbk == 32'd879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                880   :   assert (rdbk == 32'd880) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                881   :   assert (rdbk == 32'd881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                882   :   assert (rdbk == 32'd882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                883   :   assert (rdbk == 32'd883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                884   :   assert (rdbk == 32'd884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                885   :   assert (rdbk == 32'd885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                886   :   assert (rdbk == 32'd886) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                887   :   assert (rdbk == 32'd887) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                888   :   assert (rdbk == 32'd888) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                889   :   assert (rdbk == 32'd889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                890   :   assert (rdbk == 32'd890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                891   :   assert (rdbk == 32'd891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                892   :   assert (rdbk == 32'd892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                893   :   assert (rdbk == 32'd893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                894   :   assert (rdbk == 32'd894) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                895   :   assert (rdbk == 32'd895) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                896   :   assert (rdbk == 32'd896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                897   :   assert (rdbk == 32'd897) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                898   :   assert (rdbk == 32'd898) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                899   :   assert (rdbk == 32'd899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                900   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                901   :   assert (rdbk == 32'd901) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                902   :   assert (rdbk == 32'd902) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                903   :   assert (rdbk == 32'd903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                904   :   assert (rdbk == 32'd904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                905   :   assert (rdbk == 32'd905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                906   :   assert (rdbk == 32'd906) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                907   :   assert (rdbk == 32'd907) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                908   :   assert (rdbk == 32'd908) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                909   :   assert (rdbk == 32'd909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                910   :   assert (rdbk == 32'd910) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                911   :   assert (rdbk == 32'd911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                912   :   assert (rdbk == 32'd912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                913   :   assert (rdbk == 32'd913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                914   :   assert (rdbk == 32'd914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                915   :   assert (rdbk == 32'd915) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                916   :   assert (rdbk == 32'd916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                917   :   assert (rdbk == 32'd917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                918   :   assert (rdbk == 32'd918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                919   :   assert (rdbk == 32'd919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                920   :   assert (rdbk == 32'd920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                921   :   assert (rdbk == 32'd921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                922   :   assert (rdbk == 32'd922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                923   :   assert (rdbk == 32'd923) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                924   :   assert (rdbk == 32'd924) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                925   :   assert (rdbk == 32'd925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                926   :   assert (rdbk == 32'd926) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                927   :   assert (rdbk == 32'd927) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                928   :   assert (rdbk == 32'd928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                929   :   assert (rdbk == 32'd929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                930   :   assert (rdbk == 32'd930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                931   :   assert (rdbk == 32'd931) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                932   :   assert (rdbk == 32'd932) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                933   :   assert (rdbk == 32'd933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                934   :   assert (rdbk == 32'd934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                935   :   assert (rdbk == 32'd935) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                936   :   assert (rdbk == 32'd936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                937   :   assert (rdbk == 32'd937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                938   :   assert (rdbk == 32'd938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                939   :   assert (rdbk == 32'd939) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                940   :   assert (rdbk == 32'd940) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                941   :   assert (rdbk == 32'd941) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                942   :   assert (rdbk == 32'd942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                943   :   assert (rdbk == 32'd943) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                944   :   assert (rdbk == 32'd944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                945   :   assert (rdbk == 32'd945) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                946   :   assert (rdbk == 32'd946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                947   :   assert (rdbk == 32'd947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                948   :   assert (rdbk == 32'd948) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                949   :   assert (rdbk == 32'd949) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                950   :   assert (rdbk == 32'd950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                951   :   assert (rdbk == 32'd951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                952   :   assert (rdbk == 32'd952) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                953   :   assert (rdbk == 32'd953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                954   :   assert (rdbk == 32'd954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                955   :   assert (rdbk == 32'd955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                956   :   assert (rdbk == 32'd956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                957   :   assert (rdbk == 32'd957) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                958   :   assert (rdbk == 32'd958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                959   :   assert (rdbk == 32'd959) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                960   :   assert (rdbk == 32'd960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                961   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                962   :   assert (rdbk == 32'd962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                963   :   assert (rdbk == 32'd963) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                964   :   assert (rdbk == 32'd964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                965   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                966   :   assert (rdbk == 32'd966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                967   :   assert (rdbk == 32'd967) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                968   :   assert (rdbk == 32'd968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                969   :   assert (rdbk == 32'd969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                970   :   assert (rdbk == 32'd970) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                971   :   assert (rdbk == 32'd971) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                972   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                973   :   assert (rdbk == 32'd973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                974   :   assert (rdbk == 32'd974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                975   :   assert (rdbk == 32'd975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                976   :   assert (rdbk == 32'd976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                977   :   assert (rdbk == 32'd977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                978   :   assert (rdbk == 32'd978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                979   :   assert (rdbk == 32'd979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                980   :   assert (rdbk == 32'd980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                981   :   assert (rdbk == 32'd981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                982   :   assert (rdbk == 32'd982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                983   :   assert (rdbk == 32'd983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                984   :   assert (rdbk == 32'd984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                985   :   assert (rdbk == 32'd985) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                986   :   assert (rdbk == 32'd986) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                987   :   assert (rdbk == 32'd987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                988   :   assert (rdbk == 32'd988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                989   :   assert (rdbk == 32'd989) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                990   :   assert (rdbk == 32'd990) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                991   :   assert (rdbk == 32'd991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                992   :   assert (rdbk == 32'd992) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                993   :   assert (rdbk == 32'd993) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                994   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                995   :   assert (rdbk == 32'd995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                996   :   assert (rdbk == 32'd996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                997   :   assert (rdbk == 32'd997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                998   :   assert (rdbk == 32'd998) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                999   :   assert (rdbk == 32'd999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1000   :   assert (rdbk == 32'd1000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1001   :   assert (rdbk == 32'd1001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1002   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1003   :   assert (rdbk == 32'd1003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1004   :   assert (rdbk == 32'd1004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1005   :   assert (rdbk == 32'd1005) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1006   :   assert (rdbk == 32'd1006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1007   :   assert (rdbk == 32'd1007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1008   :   assert (rdbk == 32'd1008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1009   :   assert (rdbk == 32'd1009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1010   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1011   :   assert (rdbk == 32'd1011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1012   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1013   :   assert (rdbk == 32'd1013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1014   :   assert (rdbk == 32'd1014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1015   :   assert (rdbk == 32'd1015) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1016   :   assert (rdbk == 32'd1016) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1017   :   assert (rdbk == 32'd1017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1018   :   assert (rdbk == 32'd1018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1019   :   assert (rdbk == 32'd1019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1020   :   assert (rdbk == 32'd1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1021   :   assert (rdbk == 32'd1021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1022   :   assert (rdbk == 32'd1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1023   :   assert (rdbk == 32'd1023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end



        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- Pointwise-Multiplication (Dilithium)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_mul_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_mul_dilithium.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_dilithium_pointwise_mul = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+128), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd1089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd1156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd1521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd1600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd1764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd1849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd2025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd2116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd2209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd2304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd2401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd2500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd2601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd2704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd2916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd3025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd3136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd3249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd3364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd3481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd3600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd3721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd3844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd3969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd4096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd4225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd4356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd4489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd4761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd4900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd5041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd5329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd5476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd5625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd5776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd5929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd6084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd6241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd6400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd6561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd6724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd6889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd7056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd7225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd7396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd7569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd7744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd7921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd8100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd8281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd8464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd8649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd8836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd9025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd9216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd9409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd9604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd9801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd10201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd10404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd11025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd11236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd11449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd11881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd12100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd12321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd12544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd12769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd12996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd13225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd13456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd13689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd13924) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd14161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd14400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd14641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd14884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd15129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd15376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd15625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd15876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd16129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd16384) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd16641) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd16900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd17161) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd17424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd17689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd17956) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd18225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd18496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd18769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd19044) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd19321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd19600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd19881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd20164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd20449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd20736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd21025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd21316) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd21609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd21904) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd22201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd22500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd22801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd23104) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd23409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd23716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd24025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd24336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd24649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd24964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd25281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd25600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd25921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd26244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd26569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd26896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd27225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd27556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd27889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd28224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd28561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd28900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd29241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd29584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd29929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd30276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd30625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd30976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd31329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd31684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd32041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd32400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd32761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd33124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd33489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd33856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd34225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd34596) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd34969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd35344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd35721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd36100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd36481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd36864) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd37249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd37636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd38025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd38416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd38809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd39204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd39601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd40000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd40401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd40804) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd41209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd41616) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd42025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd42436) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd42849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd43264) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd43681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd44100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd44521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd44944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd45369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd45796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd46225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd46656) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd47089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd47524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd47961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd48400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd48841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd49284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd49729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd50176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd50625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd51076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd51529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd51984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd52441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd52900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd53361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd53824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd54289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd54756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd55225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd55696) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd56169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd56644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd57121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd57600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd58081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd58564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd59049) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd59536) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd60025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd60516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd61009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd61504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd62001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd62500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd63001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd63504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd64009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd64516) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd65025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- Basecase-Multiplication (Kyber)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_mul_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_mul_kyber.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_kyber_base_mul = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<256 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+256), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd3180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd12) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd2461) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd40) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd1236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd84) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd2795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd1739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd62) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd1929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd2988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd852) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd2435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd1200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd553) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd1404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd1624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd2422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd1860) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd756) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd2112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd2882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd2380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd319) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd2664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd2964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd3280) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd633) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1043) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd631) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd85) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd3155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd1375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd254) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd1771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd2527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd2611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd1624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd3055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd1157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd2638) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd1154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd1973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd1662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd2973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd2186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd1937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd2726) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd1380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd3282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd1113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd3234) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd1717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd3072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd2337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd349) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd2973) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd2850) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd2335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd1648) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd2063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd2348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd3064) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd1920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd467) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd1215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd2443) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd1979) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd1163) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd2759) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd1233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd2969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd1038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd1866) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd2710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd1267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd1117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd1086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd2009) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd3132) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd2917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd2972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd3269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd1452) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd3310) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd2408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd1718) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd51) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd1039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd2043) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd61) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd3063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd1845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd770) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd3011) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd1822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd2410) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd2890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd645) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd960) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd1745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd3105) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd2861) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd2030) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd2065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd1812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd2976) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd2608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd827) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd2023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd1627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd3235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd2799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd1134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd1418) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd2378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd2187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd1585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd2877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd3007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd856) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd2750) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd2180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd1006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd191) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd1428) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd1547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd2031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd2919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd2849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd2382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd1951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd1909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd1381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd2608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd1500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd2168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd2984) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd2942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd1155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd1250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd2671) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd2395) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd2422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd3055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd2003) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd2237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd2845) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd2010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd2116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd2110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd415) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd2188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd2059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd2357) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd390) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd414) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd2066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd1988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd2735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd2137) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd2117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd2563) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd2272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd1249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd699) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd2099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd2471) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd3297) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd930) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd2698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd2734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd3273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd1916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd3061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd1584) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd1794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd2235) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd2007) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd2695) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd1440) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd2494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd3064) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd1097) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd2309) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd3045) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd2760) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd1680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd560) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd331) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd785) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd2327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd1775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd1761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd3038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end

        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- Pointwise-Multiplication (Falcon-512)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_mul_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_mul_falcon512.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon512_pointwise_mul = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<512 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+128), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd1089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd1156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd1521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd1600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd1764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd1849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd2025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd2116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd2209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd2304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd2401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd2500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd2601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd2704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd2916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd3025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd3136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd3249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd3364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd3481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd3600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd3721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd3844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd3969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd4096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd4225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd4356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd4489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd4761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd4900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd5041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd5329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd5476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd5625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd5776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd5929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd6084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd6241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd6400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd6561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd6724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd6889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd7056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd7225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd7396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd7569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd7744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd7921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd8100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd8281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd8464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd8649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd8836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd9025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd9216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd9409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd9604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd9801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd10201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd10404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd11025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd11236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd11449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd11881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd12100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd1167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd1400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd1635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd1872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd2111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd2352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd2595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd2840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd3087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd3336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd3587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd3840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd4095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd4611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd4872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd5135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd5400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd5667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd5936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd6207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd6480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd6755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd7032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd7311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd7592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd7875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd8160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd8447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd8736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd9027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd9320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd9615) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd9912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd10211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd10512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd10815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd11120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd11427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd11736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd12047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd1343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd1991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd2318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd2647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd2978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd3311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd3646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd3983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd4322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd4663) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd5006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd5351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd5698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd6047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd6398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd6751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd7106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd7463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd7822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd8183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd8546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd8911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd9278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd9647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd10018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd10391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd10766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd11143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd11903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd12286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd1158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd1549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd1942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd2337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd2734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd3133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd3534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd3937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd4342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd4749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd5158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd5569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd5982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd6397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd6814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd7233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd7654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd8077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd8502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd8929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd9358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd10222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd10657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd11094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd11533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd11974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd1469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd1920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd2373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd2828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd3285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd3744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd4205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd4668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd5133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd5600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd6069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd6540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd7013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd7488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd7965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd8444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd8925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd9408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd9893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd10380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd10869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd11360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd11853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd1055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd1556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd2059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd2564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd3071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd3580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd4091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd4604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd5119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd5636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd6155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd6676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd7199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd7724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd8251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd8780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd9311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd9844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd10379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd10916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd11455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd11996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd1342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd1891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd2442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd2995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd3550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd4107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd4666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd5227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd5790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd6355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd6922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd7491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd8062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd8635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd9210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd9787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd10366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd10947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd11530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd12115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd1593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd2186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd2781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd3378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd3977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd4578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd5181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd5786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd6393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd7002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd7613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd8226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd8841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd9458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd10077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd10698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd11321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd11946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd1544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd2177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd2812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd3449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd4088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd4729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd5372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd6017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd6664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd7313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd7964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd8617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd9272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd9929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd10588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd11249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd11912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd1624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd2295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd2968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd3643) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd4320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd4999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd5680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd6363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd7048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd7735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd8424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd9115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd9808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd10503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd11200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd11899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd1014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd1719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd2426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd3135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd3846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd4559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd5274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd5991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd6710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd7431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd8154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd8879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd9606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd10335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd11066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd11799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd1721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd2462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd3205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd3950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd4697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd5446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd6197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd6950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd7705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd8462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd9221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd9982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd10745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd11510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd12277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd1528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd2301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd3076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd3853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd4632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd5413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd6196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd6981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd7768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd8557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd9348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd10141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd10936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd11733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd1044) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd1847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd2652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd3459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd4268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd5079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd5892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd6707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd7524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd8343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd9164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd9987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd10812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd11639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd1843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd2678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd3515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd4354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd5195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd6038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd6883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd7730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd8579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd9430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd10283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd11138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd11995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd1426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd2289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd3154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd4021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd4890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd5761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd6634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd7509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd8386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd9265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd10146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd11029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd11914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd1401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd2292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd3185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd4080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd4977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd5876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd6777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd7680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd8585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd9492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd10401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd11312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd12225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd1768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd2687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd3608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd4531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd5456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd6383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd7312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd8243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd9176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd10111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd11048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd11987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd1582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd2527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd3474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd4423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd5374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd6327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd7282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd8239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd9198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd10159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd11122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd12087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd1734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd2705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd3678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd4653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd5630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd6609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd7590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd8573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd9558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd10545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd11534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd1229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd2224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd3221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd4220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd5221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd6224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd7229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd8236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd9245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd10256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd11269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd12284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd2031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd3052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end


        $fwrite(f,"----------------------------------------------------------------\n");   
        $fwrite(f,"-- Pointwise-Multiplication (Falcon-1024)\n");
        $fwrite(f,"----------------------------------------------------------------\n");   
             
        // Write IMEM from File
        write_imem_from_file_tl_ul(.log_filehandle(f), .imem_file_path({mem_path, "imem_mul_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        $fwrite(f,"-- IMEM\n");
        // Read IMEM  
        for (int i=0 ; i<129 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_IMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end     
 
         // Write DMEM from File
        write_dmem_from_file_tl_ul(.log_filehandle(f), .dmem_file_path({mem_path, "dmem_mul_falcon1024.txt"}), .clk(clk_i), .clk_cycles(cc), .start_address(0), .tl_o(tl_o), .tl_i(tl_i_d) );

        $fwrite(f,"-- DMEM\n");
        // Read DMEM  
        for (int i=0 ; i<16 ; i++) begin 
            //read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i), .tl_o(tl_o), .tl_i(tl_i_d) );
        end   
                   
        $fwrite(f,"----------------------------------------------------------------\n");   
  
        // Set Instruction Counter to zero (optional)
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h0), .address(OTBN_INSN_CNT_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        
        // Start Programm in IMEM
        write_tl_ul(.log_filehandle(f), .clk(clk_i), .clk_cycles(cc), .data(32'h1), .address(OTBN_CMD_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        cc_start = cc;
        // Poll on Status Register until Programm is finished
        rdbk = '1;
        while (rdbk != '0) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_STATUS_OFFSET), .tl_o(tl_o), .tl_i(tl_i_d) );
        end 
        
        // Measure CC
        cc_stop = cc; 
        cc_count_falcon1024_pointwise_mul = cc_stop - cc_start;        
               
        // Read DMEM  
        for (int i=0 ; i<1024 ; i++) begin 
            read_tl_ul(.log_filehandle(f), .data(rdbk), .clk(clk_i), .clk_cycles(cc), .address(OTBN_DMEM_OFFSET+4*i+128), .tl_o(tl_o), .tl_i(tl_i_d) );
            
            case(i)
                0   :   assert (rdbk == 32'd0) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1   :   assert (rdbk == 32'd1) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                2   :   assert (rdbk == 32'd4) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                3   :   assert (rdbk == 32'd9) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                4   :   assert (rdbk == 32'd16) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                5   :   assert (rdbk == 32'd25) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                6   :   assert (rdbk == 32'd36) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                7   :   assert (rdbk == 32'd49) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                8   :   assert (rdbk == 32'd64) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                9   :   assert (rdbk == 32'd81) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                10   :   assert (rdbk == 32'd100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                11   :   assert (rdbk == 32'd121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                12   :   assert (rdbk == 32'd144) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                13   :   assert (rdbk == 32'd169) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                14   :   assert (rdbk == 32'd196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                15   :   assert (rdbk == 32'd225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                16   :   assert (rdbk == 32'd256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                17   :   assert (rdbk == 32'd289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                18   :   assert (rdbk == 32'd324) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                19   :   assert (rdbk == 32'd361) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                20   :   assert (rdbk == 32'd400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                21   :   assert (rdbk == 32'd441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                22   :   assert (rdbk == 32'd484) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                23   :   assert (rdbk == 32'd529) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                24   :   assert (rdbk == 32'd576) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                25   :   assert (rdbk == 32'd625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                26   :   assert (rdbk == 32'd676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                27   :   assert (rdbk == 32'd729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                28   :   assert (rdbk == 32'd784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                29   :   assert (rdbk == 32'd841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                30   :   assert (rdbk == 32'd900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                31   :   assert (rdbk == 32'd961) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                32   :   assert (rdbk == 32'd1024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                33   :   assert (rdbk == 32'd1089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                34   :   assert (rdbk == 32'd1156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                35   :   assert (rdbk == 32'd1225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                36   :   assert (rdbk == 32'd1296) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                37   :   assert (rdbk == 32'd1369) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                38   :   assert (rdbk == 32'd1444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                39   :   assert (rdbk == 32'd1521) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                40   :   assert (rdbk == 32'd1600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                41   :   assert (rdbk == 32'd1681) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                42   :   assert (rdbk == 32'd1764) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                43   :   assert (rdbk == 32'd1849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                44   :   assert (rdbk == 32'd1936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                45   :   assert (rdbk == 32'd2025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                46   :   assert (rdbk == 32'd2116) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                47   :   assert (rdbk == 32'd2209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                48   :   assert (rdbk == 32'd2304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                49   :   assert (rdbk == 32'd2401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                50   :   assert (rdbk == 32'd2500) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                51   :   assert (rdbk == 32'd2601) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                52   :   assert (rdbk == 32'd2704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                53   :   assert (rdbk == 32'd2809) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                54   :   assert (rdbk == 32'd2916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                55   :   assert (rdbk == 32'd3025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                56   :   assert (rdbk == 32'd3136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                57   :   assert (rdbk == 32'd3249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                58   :   assert (rdbk == 32'd3364) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                59   :   assert (rdbk == 32'd3481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                60   :   assert (rdbk == 32'd3600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                61   :   assert (rdbk == 32'd3721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                62   :   assert (rdbk == 32'd3844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                63   :   assert (rdbk == 32'd3969) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                64   :   assert (rdbk == 32'd4096) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                65   :   assert (rdbk == 32'd4225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                66   :   assert (rdbk == 32'd4356) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                67   :   assert (rdbk == 32'd4489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                68   :   assert (rdbk == 32'd4624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                69   :   assert (rdbk == 32'd4761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                70   :   assert (rdbk == 32'd4900) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                71   :   assert (rdbk == 32'd5041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                72   :   assert (rdbk == 32'd5184) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                73   :   assert (rdbk == 32'd5329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                74   :   assert (rdbk == 32'd5476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                75   :   assert (rdbk == 32'd5625) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                76   :   assert (rdbk == 32'd5776) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                77   :   assert (rdbk == 32'd5929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                78   :   assert (rdbk == 32'd6084) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                79   :   assert (rdbk == 32'd6241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                80   :   assert (rdbk == 32'd6400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                81   :   assert (rdbk == 32'd6561) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                82   :   assert (rdbk == 32'd6724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                83   :   assert (rdbk == 32'd6889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                84   :   assert (rdbk == 32'd7056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                85   :   assert (rdbk == 32'd7225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                86   :   assert (rdbk == 32'd7396) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                87   :   assert (rdbk == 32'd7569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                88   :   assert (rdbk == 32'd7744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                89   :   assert (rdbk == 32'd7921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                90   :   assert (rdbk == 32'd8100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                91   :   assert (rdbk == 32'd8281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                92   :   assert (rdbk == 32'd8464) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                93   :   assert (rdbk == 32'd8649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                94   :   assert (rdbk == 32'd8836) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                95   :   assert (rdbk == 32'd9025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                96   :   assert (rdbk == 32'd9216) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                97   :   assert (rdbk == 32'd9409) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                98   :   assert (rdbk == 32'd9604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                99   :   assert (rdbk == 32'd9801) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                100   :   assert (rdbk == 32'd10000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                101   :   assert (rdbk == 32'd10201) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                102   :   assert (rdbk == 32'd10404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                103   :   assert (rdbk == 32'd10609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                104   :   assert (rdbk == 32'd10816) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                105   :   assert (rdbk == 32'd11025) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                106   :   assert (rdbk == 32'd11236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                107   :   assert (rdbk == 32'd11449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                108   :   assert (rdbk == 32'd11664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                109   :   assert (rdbk == 32'd11881) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                110   :   assert (rdbk == 32'd12100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                111   :   assert (rdbk == 32'd32) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                112   :   assert (rdbk == 32'd255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                113   :   assert (rdbk == 32'd480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                114   :   assert (rdbk == 32'd707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                115   :   assert (rdbk == 32'd936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                116   :   assert (rdbk == 32'd1167) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                117   :   assert (rdbk == 32'd1400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                118   :   assert (rdbk == 32'd1635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                119   :   assert (rdbk == 32'd1872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                120   :   assert (rdbk == 32'd2111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                121   :   assert (rdbk == 32'd2352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                122   :   assert (rdbk == 32'd2595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                123   :   assert (rdbk == 32'd2840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                124   :   assert (rdbk == 32'd3087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                125   :   assert (rdbk == 32'd3336) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                126   :   assert (rdbk == 32'd3587) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                127   :   assert (rdbk == 32'd3840) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                128   :   assert (rdbk == 32'd4095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                129   :   assert (rdbk == 32'd4352) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                130   :   assert (rdbk == 32'd4611) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                131   :   assert (rdbk == 32'd4872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                132   :   assert (rdbk == 32'd5135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                133   :   assert (rdbk == 32'd5400) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                134   :   assert (rdbk == 32'd5667) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                135   :   assert (rdbk == 32'd5936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                136   :   assert (rdbk == 32'd6207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                137   :   assert (rdbk == 32'd6480) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                138   :   assert (rdbk == 32'd6755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                139   :   assert (rdbk == 32'd7032) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                140   :   assert (rdbk == 32'd7311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                141   :   assert (rdbk == 32'd7592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                142   :   assert (rdbk == 32'd7875) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                143   :   assert (rdbk == 32'd8160) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                144   :   assert (rdbk == 32'd8447) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                145   :   assert (rdbk == 32'd8736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                146   :   assert (rdbk == 32'd9027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                147   :   assert (rdbk == 32'd9320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                148   :   assert (rdbk == 32'd9615) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                149   :   assert (rdbk == 32'd9912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                150   :   assert (rdbk == 32'd10211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                151   :   assert (rdbk == 32'd10512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                152   :   assert (rdbk == 32'd10815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                153   :   assert (rdbk == 32'd11120) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                154   :   assert (rdbk == 32'd11427) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                155   :   assert (rdbk == 32'd11736) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                156   :   assert (rdbk == 32'd12047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                157   :   assert (rdbk == 32'd71) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                158   :   assert (rdbk == 32'd386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                159   :   assert (rdbk == 32'd703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                160   :   assert (rdbk == 32'd1022) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                161   :   assert (rdbk == 32'd1343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                162   :   assert (rdbk == 32'd1666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                163   :   assert (rdbk == 32'd1991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                164   :   assert (rdbk == 32'd2318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                165   :   assert (rdbk == 32'd2647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                166   :   assert (rdbk == 32'd2978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                167   :   assert (rdbk == 32'd3311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                168   :   assert (rdbk == 32'd3646) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                169   :   assert (rdbk == 32'd3983) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                170   :   assert (rdbk == 32'd4322) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                171   :   assert (rdbk == 32'd4663) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                172   :   assert (rdbk == 32'd5006) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                173   :   assert (rdbk == 32'd5351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                174   :   assert (rdbk == 32'd5698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                175   :   assert (rdbk == 32'd6047) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                176   :   assert (rdbk == 32'd6398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                177   :   assert (rdbk == 32'd6751) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                178   :   assert (rdbk == 32'd7106) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                179   :   assert (rdbk == 32'd7463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                180   :   assert (rdbk == 32'd7822) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                181   :   assert (rdbk == 32'd8183) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                182   :   assert (rdbk == 32'd8546) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                183   :   assert (rdbk == 32'd8911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                184   :   assert (rdbk == 32'd9278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                185   :   assert (rdbk == 32'd9647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                186   :   assert (rdbk == 32'd10018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                187   :   assert (rdbk == 32'd10391) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                188   :   assert (rdbk == 32'd10766) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                189   :   assert (rdbk == 32'd11143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                190   :   assert (rdbk == 32'd11522) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                191   :   assert (rdbk == 32'd11903) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                192   :   assert (rdbk == 32'd12286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                193   :   assert (rdbk == 32'd382) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                194   :   assert (rdbk == 32'd769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                195   :   assert (rdbk == 32'd1158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                196   :   assert (rdbk == 32'd1549) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                197   :   assert (rdbk == 32'd1942) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                198   :   assert (rdbk == 32'd2337) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                199   :   assert (rdbk == 32'd2734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                200   :   assert (rdbk == 32'd3133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                201   :   assert (rdbk == 32'd3534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                202   :   assert (rdbk == 32'd3937) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                203   :   assert (rdbk == 32'd4342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                204   :   assert (rdbk == 32'd4749) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                205   :   assert (rdbk == 32'd5158) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                206   :   assert (rdbk == 32'd5569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                207   :   assert (rdbk == 32'd5982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                208   :   assert (rdbk == 32'd6397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                209   :   assert (rdbk == 32'd6814) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                210   :   assert (rdbk == 32'd7233) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                211   :   assert (rdbk == 32'd7654) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                212   :   assert (rdbk == 32'd8077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                213   :   assert (rdbk == 32'd8502) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                214   :   assert (rdbk == 32'd8929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                215   :   assert (rdbk == 32'd9358) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                216   :   assert (rdbk == 32'd9789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                217   :   assert (rdbk == 32'd10222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                218   :   assert (rdbk == 32'd10657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                219   :   assert (rdbk == 32'd11094) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                220   :   assert (rdbk == 32'd11533) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                221   :   assert (rdbk == 32'd11974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                222   :   assert (rdbk == 32'd128) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                223   :   assert (rdbk == 32'd573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                224   :   assert (rdbk == 32'd1020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                225   :   assert (rdbk == 32'd1469) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                226   :   assert (rdbk == 32'd1920) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                227   :   assert (rdbk == 32'd2373) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                228   :   assert (rdbk == 32'd2828) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                229   :   assert (rdbk == 32'd3285) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                230   :   assert (rdbk == 32'd3744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                231   :   assert (rdbk == 32'd4205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                232   :   assert (rdbk == 32'd4668) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                233   :   assert (rdbk == 32'd5133) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                234   :   assert (rdbk == 32'd5600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                235   :   assert (rdbk == 32'd6069) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                236   :   assert (rdbk == 32'd6540) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                237   :   assert (rdbk == 32'd7013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                238   :   assert (rdbk == 32'd7488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                239   :   assert (rdbk == 32'd7965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                240   :   assert (rdbk == 32'd8444) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                241   :   assert (rdbk == 32'd8925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                242   :   assert (rdbk == 32'd9408) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                243   :   assert (rdbk == 32'd9893) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                244   :   assert (rdbk == 32'd10380) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                245   :   assert (rdbk == 32'd10869) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                246   :   assert (rdbk == 32'd11360) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                247   :   assert (rdbk == 32'd11853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                248   :   assert (rdbk == 32'd59) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                249   :   assert (rdbk == 32'd556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                250   :   assert (rdbk == 32'd1055) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                251   :   assert (rdbk == 32'd1556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                252   :   assert (rdbk == 32'd2059) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                253   :   assert (rdbk == 32'd2564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                254   :   assert (rdbk == 32'd3071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                255   :   assert (rdbk == 32'd3580) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                256   :   assert (rdbk == 32'd4091) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                257   :   assert (rdbk == 32'd4604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                258   :   assert (rdbk == 32'd5119) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                259   :   assert (rdbk == 32'd5636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                260   :   assert (rdbk == 32'd6155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                261   :   assert (rdbk == 32'd6676) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                262   :   assert (rdbk == 32'd7199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                263   :   assert (rdbk == 32'd7724) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                264   :   assert (rdbk == 32'd8251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                265   :   assert (rdbk == 32'd8780) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                266   :   assert (rdbk == 32'd9311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                267   :   assert (rdbk == 32'd9844) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                268   :   assert (rdbk == 32'd10379) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                269   :   assert (rdbk == 32'd10916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                270   :   assert (rdbk == 32'd11455) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                271   :   assert (rdbk == 32'd11996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                272   :   assert (rdbk == 32'd250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                273   :   assert (rdbk == 32'd795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                274   :   assert (rdbk == 32'd1342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                275   :   assert (rdbk == 32'd1891) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                276   :   assert (rdbk == 32'd2442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                277   :   assert (rdbk == 32'd2995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                278   :   assert (rdbk == 32'd3550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                279   :   assert (rdbk == 32'd4107) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                280   :   assert (rdbk == 32'd4666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                281   :   assert (rdbk == 32'd5227) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                282   :   assert (rdbk == 32'd5790) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                283   :   assert (rdbk == 32'd6355) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                284   :   assert (rdbk == 32'd6922) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                285   :   assert (rdbk == 32'd7491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                286   :   assert (rdbk == 32'd8062) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                287   :   assert (rdbk == 32'd8635) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                288   :   assert (rdbk == 32'd9210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                289   :   assert (rdbk == 32'd9787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                290   :   assert (rdbk == 32'd10366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                291   :   assert (rdbk == 32'd10947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                292   :   assert (rdbk == 32'd11530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                293   :   assert (rdbk == 32'd12115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                294   :   assert (rdbk == 32'd413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                295   :   assert (rdbk == 32'd1002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                296   :   assert (rdbk == 32'd1593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                297   :   assert (rdbk == 32'd2186) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                298   :   assert (rdbk == 32'd2781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                299   :   assert (rdbk == 32'd3378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                300   :   assert (rdbk == 32'd3977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                301   :   assert (rdbk == 32'd4578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                302   :   assert (rdbk == 32'd5181) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                303   :   assert (rdbk == 32'd5786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                304   :   assert (rdbk == 32'd6393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                305   :   assert (rdbk == 32'd7002) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                306   :   assert (rdbk == 32'd7613) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                307   :   assert (rdbk == 32'd8226) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                308   :   assert (rdbk == 32'd8841) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                309   :   assert (rdbk == 32'd9458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                310   :   assert (rdbk == 32'd10077) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                311   :   assert (rdbk == 32'd10698) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                312   :   assert (rdbk == 32'd11321) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                313   :   assert (rdbk == 32'd11946) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                314   :   assert (rdbk == 32'd284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                315   :   assert (rdbk == 32'd913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                316   :   assert (rdbk == 32'd1544) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                317   :   assert (rdbk == 32'd2177) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                318   :   assert (rdbk == 32'd2812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                319   :   assert (rdbk == 32'd3449) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                320   :   assert (rdbk == 32'd4088) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                321   :   assert (rdbk == 32'd4729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                322   :   assert (rdbk == 32'd5372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                323   :   assert (rdbk == 32'd6017) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                324   :   assert (rdbk == 32'd6664) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                325   :   assert (rdbk == 32'd7313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                326   :   assert (rdbk == 32'd7964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                327   :   assert (rdbk == 32'd8617) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                328   :   assert (rdbk == 32'd9272) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                329   :   assert (rdbk == 32'd9929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                330   :   assert (rdbk == 32'd10588) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                331   :   assert (rdbk == 32'd11249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                332   :   assert (rdbk == 32'd11912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                333   :   assert (rdbk == 32'd288) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                334   :   assert (rdbk == 32'd955) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                335   :   assert (rdbk == 32'd1624) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                336   :   assert (rdbk == 32'd2295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                337   :   assert (rdbk == 32'd2968) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                338   :   assert (rdbk == 32'd3643) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                339   :   assert (rdbk == 32'd4320) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                340   :   assert (rdbk == 32'd4999) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                341   :   assert (rdbk == 32'd5680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                342   :   assert (rdbk == 32'd6363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                343   :   assert (rdbk == 32'd7048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                344   :   assert (rdbk == 32'd7735) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                345   :   assert (rdbk == 32'd8424) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                346   :   assert (rdbk == 32'd9115) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                347   :   assert (rdbk == 32'd9808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                348   :   assert (rdbk == 32'd10503) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                349   :   assert (rdbk == 32'd11200) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                350   :   assert (rdbk == 32'd11899) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                351   :   assert (rdbk == 32'd311) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                352   :   assert (rdbk == 32'd1014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                353   :   assert (rdbk == 32'd1719) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                354   :   assert (rdbk == 32'd2426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                355   :   assert (rdbk == 32'd3135) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                356   :   assert (rdbk == 32'd3846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                357   :   assert (rdbk == 32'd4559) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                358   :   assert (rdbk == 32'd5274) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                359   :   assert (rdbk == 32'd5991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                360   :   assert (rdbk == 32'd6710) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                361   :   assert (rdbk == 32'd7431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                362   :   assert (rdbk == 32'd8154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                363   :   assert (rdbk == 32'd8879) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                364   :   assert (rdbk == 32'd9606) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                365   :   assert (rdbk == 32'd10335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                366   :   assert (rdbk == 32'd11066) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                367   :   assert (rdbk == 32'd11799) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                368   :   assert (rdbk == 32'd245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                369   :   assert (rdbk == 32'd982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                370   :   assert (rdbk == 32'd1721) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                371   :   assert (rdbk == 32'd2462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                372   :   assert (rdbk == 32'd3205) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                373   :   assert (rdbk == 32'd3950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                374   :   assert (rdbk == 32'd4697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                375   :   assert (rdbk == 32'd5446) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                376   :   assert (rdbk == 32'd6197) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                377   :   assert (rdbk == 32'd6950) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                378   :   assert (rdbk == 32'd7705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                379   :   assert (rdbk == 32'd8462) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                380   :   assert (rdbk == 32'd9221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                381   :   assert (rdbk == 32'd9982) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                382   :   assert (rdbk == 32'd10745) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                383   :   assert (rdbk == 32'd11510) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                384   :   assert (rdbk == 32'd12277) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                385   :   assert (rdbk == 32'd757) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                386   :   assert (rdbk == 32'd1528) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                387   :   assert (rdbk == 32'd2301) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                388   :   assert (rdbk == 32'd3076) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                389   :   assert (rdbk == 32'd3853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                390   :   assert (rdbk == 32'd4632) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                391   :   assert (rdbk == 32'd5413) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                392   :   assert (rdbk == 32'd6196) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                393   :   assert (rdbk == 32'd6981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                394   :   assert (rdbk == 32'd7768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                395   :   assert (rdbk == 32'd8557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                396   :   assert (rdbk == 32'd9348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                397   :   assert (rdbk == 32'd10141) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                398   :   assert (rdbk == 32'd10936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                399   :   assert (rdbk == 32'd11733) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                400   :   assert (rdbk == 32'd243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                401   :   assert (rdbk == 32'd1044) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                402   :   assert (rdbk == 32'd1847) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                403   :   assert (rdbk == 32'd2652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                404   :   assert (rdbk == 32'd3459) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                405   :   assert (rdbk == 32'd4268) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                406   :   assert (rdbk == 32'd5079) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                407   :   assert (rdbk == 32'd5892) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                408   :   assert (rdbk == 32'd6707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                409   :   assert (rdbk == 32'd7524) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                410   :   assert (rdbk == 32'd8343) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                411   :   assert (rdbk == 32'd9164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                412   :   assert (rdbk == 32'd9987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                413   :   assert (rdbk == 32'd10812) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                414   :   assert (rdbk == 32'd11639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                415   :   assert (rdbk == 32'd179) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                416   :   assert (rdbk == 32'd1010) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                417   :   assert (rdbk == 32'd1843) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                418   :   assert (rdbk == 32'd2678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                419   :   assert (rdbk == 32'd3515) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                420   :   assert (rdbk == 32'd4354) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                421   :   assert (rdbk == 32'd5195) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                422   :   assert (rdbk == 32'd6038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                423   :   assert (rdbk == 32'd6883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                424   :   assert (rdbk == 32'd7730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                425   :   assert (rdbk == 32'd8579) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                426   :   assert (rdbk == 32'd9430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                427   :   assert (rdbk == 32'd10283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                428   :   assert (rdbk == 32'd11138) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                429   :   assert (rdbk == 32'd11995) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                430   :   assert (rdbk == 32'd565) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                431   :   assert (rdbk == 32'd1426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                432   :   assert (rdbk == 32'd2289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                433   :   assert (rdbk == 32'd3154) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                434   :   assert (rdbk == 32'd4021) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                435   :   assert (rdbk == 32'd4890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                436   :   assert (rdbk == 32'd5761) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                437   :   assert (rdbk == 32'd6634) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                438   :   assert (rdbk == 32'd7509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                439   :   assert (rdbk == 32'd8386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                440   :   assert (rdbk == 32'd9265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                441   :   assert (rdbk == 32'd10146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                442   :   assert (rdbk == 32'd11029) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                443   :   assert (rdbk == 32'd11914) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                444   :   assert (rdbk == 32'd512) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                445   :   assert (rdbk == 32'd1401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                446   :   assert (rdbk == 32'd2292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                447   :   assert (rdbk == 32'd3185) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                448   :   assert (rdbk == 32'd4080) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                449   :   assert (rdbk == 32'd4977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                450   :   assert (rdbk == 32'd5876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                451   :   assert (rdbk == 32'd6777) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                452   :   assert (rdbk == 32'd7680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                453   :   assert (rdbk == 32'd8585) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                454   :   assert (rdbk == 32'd9492) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                455   :   assert (rdbk == 32'd10401) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                456   :   assert (rdbk == 32'd11312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                457   :   assert (rdbk == 32'd12225) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                458   :   assert (rdbk == 32'd851) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                459   :   assert (rdbk == 32'd1768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                460   :   assert (rdbk == 32'd2687) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                461   :   assert (rdbk == 32'd3608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                462   :   assert (rdbk == 32'd4531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                463   :   assert (rdbk == 32'd5456) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                464   :   assert (rdbk == 32'd6383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                465   :   assert (rdbk == 32'd7312) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                466   :   assert (rdbk == 32'd8243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                467   :   assert (rdbk == 32'd9176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                468   :   assert (rdbk == 32'd10111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                469   :   assert (rdbk == 32'd11048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                470   :   assert (rdbk == 32'd11987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                471   :   assert (rdbk == 32'd639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                472   :   assert (rdbk == 32'd1582) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                473   :   assert (rdbk == 32'd2527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                474   :   assert (rdbk == 32'd3474) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                475   :   assert (rdbk == 32'd4423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                476   :   assert (rdbk == 32'd5374) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                477   :   assert (rdbk == 32'd6327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                478   :   assert (rdbk == 32'd7282) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                479   :   assert (rdbk == 32'd8239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                480   :   assert (rdbk == 32'd9198) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                481   :   assert (rdbk == 32'd10159) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                482   :   assert (rdbk == 32'd11122) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                483   :   assert (rdbk == 32'd12087) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                484   :   assert (rdbk == 32'd765) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                485   :   assert (rdbk == 32'd1734) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                486   :   assert (rdbk == 32'd2705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                487   :   assert (rdbk == 32'd3678) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                488   :   assert (rdbk == 32'd4653) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                489   :   assert (rdbk == 32'd5630) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                490   :   assert (rdbk == 32'd6609) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                491   :   assert (rdbk == 32'd7590) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                492   :   assert (rdbk == 32'd8573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                493   :   assert (rdbk == 32'd9558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                494   :   assert (rdbk == 32'd10545) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                495   :   assert (rdbk == 32'd11534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                496   :   assert (rdbk == 32'd236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                497   :   assert (rdbk == 32'd1229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                498   :   assert (rdbk == 32'd2224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                499   :   assert (rdbk == 32'd3221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                500   :   assert (rdbk == 32'd4220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                501   :   assert (rdbk == 32'd5221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                502   :   assert (rdbk == 32'd6224) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                503   :   assert (rdbk == 32'd7229) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                504   :   assert (rdbk == 32'd8236) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                505   :   assert (rdbk == 32'd9245) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                506   :   assert (rdbk == 32'd10256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                507   :   assert (rdbk == 32'd11269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                508   :   assert (rdbk == 32'd12284) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                509   :   assert (rdbk == 32'd1012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                510   :   assert (rdbk == 32'd2031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                511   :   assert (rdbk == 32'd3052) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                512   :   assert (rdbk == 32'd4075) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                513   :   assert (rdbk == 32'd5100) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                514   :   assert (rdbk == 32'd6127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                515   :   assert (rdbk == 32'd7156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                516   :   assert (rdbk == 32'd8187) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                517   :   assert (rdbk == 32'd9220) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                518   :   assert (rdbk == 32'd10255) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                519   :   assert (rdbk == 32'd11292) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                520   :   assert (rdbk == 32'd42) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                521   :   assert (rdbk == 32'd1083) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                522   :   assert (rdbk == 32'd2126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                523   :   assert (rdbk == 32'd3171) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                524   :   assert (rdbk == 32'd4218) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                525   :   assert (rdbk == 32'd5267) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                526   :   assert (rdbk == 32'd6318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                527   :   assert (rdbk == 32'd7371) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                528   :   assert (rdbk == 32'd8426) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                529   :   assert (rdbk == 32'd9483) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                530   :   assert (rdbk == 32'd10542) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                531   :   assert (rdbk == 32'd11603) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                532   :   assert (rdbk == 32'd377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                533   :   assert (rdbk == 32'd1442) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                534   :   assert (rdbk == 32'd2509) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                535   :   assert (rdbk == 32'd3578) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                536   :   assert (rdbk == 32'd4649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                537   :   assert (rdbk == 32'd5722) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                538   :   assert (rdbk == 32'd6797) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                539   :   assert (rdbk == 32'd7874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                540   :   assert (rdbk == 32'd8953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                541   :   assert (rdbk == 32'd10034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                542   :   assert (rdbk == 32'd11117) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                543   :   assert (rdbk == 32'd12202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                544   :   assert (rdbk == 32'd1000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                545   :   assert (rdbk == 32'd2089) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                546   :   assert (rdbk == 32'd3180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                547   :   assert (rdbk == 32'd4273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                548   :   assert (rdbk == 32'd5368) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                549   :   assert (rdbk == 32'd6465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                550   :   assert (rdbk == 32'd7564) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                551   :   assert (rdbk == 32'd8665) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                552   :   assert (rdbk == 32'd9768) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                553   :   assert (rdbk == 32'd10873) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                554   :   assert (rdbk == 32'd11980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                555   :   assert (rdbk == 32'd800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                556   :   assert (rdbk == 32'd1911) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                557   :   assert (rdbk == 32'd3024) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                558   :   assert (rdbk == 32'd4139) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                559   :   assert (rdbk == 32'd5256) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                560   :   assert (rdbk == 32'd6375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                561   :   assert (rdbk == 32'd7496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                562   :   assert (rdbk == 32'd8619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                563   :   assert (rdbk == 32'd9744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                564   :   assert (rdbk == 32'd10871) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                565   :   assert (rdbk == 32'd12000) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                566   :   assert (rdbk == 32'd842) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                567   :   assert (rdbk == 32'd1975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                568   :   assert (rdbk == 32'd3110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                569   :   assert (rdbk == 32'd4247) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                570   :   assert (rdbk == 32'd5386) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                571   :   assert (rdbk == 32'd6527) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                572   :   assert (rdbk == 32'd7670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                573   :   assert (rdbk == 32'd8815) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                574   :   assert (rdbk == 32'd9962) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                575   :   assert (rdbk == 32'd11111) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                576   :   assert (rdbk == 32'd12262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                577   :   assert (rdbk == 32'd1126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                578   :   assert (rdbk == 32'd2281) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                579   :   assert (rdbk == 32'd3438) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                580   :   assert (rdbk == 32'd4597) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                581   :   assert (rdbk == 32'd5758) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                582   :   assert (rdbk == 32'd6921) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                583   :   assert (rdbk == 32'd8086) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                584   :   assert (rdbk == 32'd9253) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                585   :   assert (rdbk == 32'd10422) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                586   :   assert (rdbk == 32'd11593) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                587   :   assert (rdbk == 32'd477) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                588   :   assert (rdbk == 32'd1652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                589   :   assert (rdbk == 32'd2829) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                590   :   assert (rdbk == 32'd4008) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                591   :   assert (rdbk == 32'd5189) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                592   :   assert (rdbk == 32'd6372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                593   :   assert (rdbk == 32'd7557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                594   :   assert (rdbk == 32'd8744) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                595   :   assert (rdbk == 32'd9933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                596   :   assert (rdbk == 32'd11124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                597   :   assert (rdbk == 32'd28) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                598   :   assert (rdbk == 32'd1223) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                599   :   assert (rdbk == 32'd2420) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                600   :   assert (rdbk == 32'd3619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                601   :   assert (rdbk == 32'd4820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                602   :   assert (rdbk == 32'd6023) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                603   :   assert (rdbk == 32'd7228) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                604   :   assert (rdbk == 32'd8435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                605   :   assert (rdbk == 32'd9644) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                606   :   assert (rdbk == 32'd10855) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                607   :   assert (rdbk == 32'd12068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                608   :   assert (rdbk == 32'd994) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                609   :   assert (rdbk == 32'd2211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                610   :   assert (rdbk == 32'd3430) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                611   :   assert (rdbk == 32'd4651) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                612   :   assert (rdbk == 32'd5874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                613   :   assert (rdbk == 32'd7099) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                614   :   assert (rdbk == 32'd8326) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                615   :   assert (rdbk == 32'd9555) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                616   :   assert (rdbk == 32'd10786) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                617   :   assert (rdbk == 32'd12019) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                618   :   assert (rdbk == 32'd965) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                619   :   assert (rdbk == 32'd2202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                620   :   assert (rdbk == 32'd3441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                621   :   assert (rdbk == 32'd4682) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                622   :   assert (rdbk == 32'd5925) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                623   :   assert (rdbk == 32'd7170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                624   :   assert (rdbk == 32'd8417) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                625   :   assert (rdbk == 32'd9666) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                626   :   assert (rdbk == 32'd10917) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                627   :   assert (rdbk == 32'd12170) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                628   :   assert (rdbk == 32'd1136) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                629   :   assert (rdbk == 32'd2393) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                630   :   assert (rdbk == 32'd3652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                631   :   assert (rdbk == 32'd4913) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                632   :   assert (rdbk == 32'd6176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                633   :   assert (rdbk == 32'd7441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                634   :   assert (rdbk == 32'd8708) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                635   :   assert (rdbk == 32'd9977) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                636   :   assert (rdbk == 32'd11248) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                637   :   assert (rdbk == 32'd232) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                638   :   assert (rdbk == 32'd1507) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                639   :   assert (rdbk == 32'd2784) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                640   :   assert (rdbk == 32'd4063) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                641   :   assert (rdbk == 32'd5344) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                642   :   assert (rdbk == 32'd6627) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                643   :   assert (rdbk == 32'd7912) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                644   :   assert (rdbk == 32'd9199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                645   :   assert (rdbk == 32'd10488) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                646   :   assert (rdbk == 32'd11779) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                647   :   assert (rdbk == 32'd783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                648   :   assert (rdbk == 32'd2078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                649   :   assert (rdbk == 32'd3375) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                650   :   assert (rdbk == 32'd4674) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                651   :   assert (rdbk == 32'd5975) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                652   :   assert (rdbk == 32'd7278) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                653   :   assert (rdbk == 32'd8583) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                654   :   assert (rdbk == 32'd9890) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                655   :   assert (rdbk == 32'd11199) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                656   :   assert (rdbk == 32'd221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                657   :   assert (rdbk == 32'd1534) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                658   :   assert (rdbk == 32'd2849) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                659   :   assert (rdbk == 32'd4166) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                660   :   assert (rdbk == 32'd5485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                661   :   assert (rdbk == 32'd6806) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                662   :   assert (rdbk == 32'd8129) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                663   :   assert (rdbk == 32'd9454) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                664   :   assert (rdbk == 32'd10781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                665   :   assert (rdbk == 32'd12110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                666   :   assert (rdbk == 32'd1152) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                667   :   assert (rdbk == 32'd2485) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                668   :   assert (rdbk == 32'd3820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                669   :   assert (rdbk == 32'd5157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                670   :   assert (rdbk == 32'd6496) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                671   :   assert (rdbk == 32'd7837) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                672   :   assert (rdbk == 32'd9180) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                673   :   assert (rdbk == 32'd10525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                674   :   assert (rdbk == 32'd11872) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                675   :   assert (rdbk == 32'd932) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                676   :   assert (rdbk == 32'd2283) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                677   :   assert (rdbk == 32'd3636) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                678   :   assert (rdbk == 32'd4991) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                679   :   assert (rdbk == 32'd6348) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                680   :   assert (rdbk == 32'd7707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                681   :   assert (rdbk == 32'd9068) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                682   :   assert (rdbk == 32'd10431) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                683   :   assert (rdbk == 32'd11796) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                684   :   assert (rdbk == 32'd874) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                685   :   assert (rdbk == 32'd2243) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                686   :   assert (rdbk == 32'd3614) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                687   :   assert (rdbk == 32'd4987) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                688   :   assert (rdbk == 32'd6362) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                689   :   assert (rdbk == 32'd7739) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                690   :   assert (rdbk == 32'd9118) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                691   :   assert (rdbk == 32'd10499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                692   :   assert (rdbk == 32'd11882) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                693   :   assert (rdbk == 32'd978) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                694   :   assert (rdbk == 32'd2365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                695   :   assert (rdbk == 32'd3754) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                696   :   assert (rdbk == 32'd5145) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                697   :   assert (rdbk == 32'd6538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                698   :   assert (rdbk == 32'd7933) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                699   :   assert (rdbk == 32'd9330) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                700   :   assert (rdbk == 32'd10729) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                701   :   assert (rdbk == 32'd12130) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                702   :   assert (rdbk == 32'd1244) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                703   :   assert (rdbk == 32'd2649) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                704   :   assert (rdbk == 32'd4056) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                705   :   assert (rdbk == 32'd5465) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                706   :   assert (rdbk == 32'd6876) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                707   :   assert (rdbk == 32'd8289) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                708   :   assert (rdbk == 32'd9704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                709   :   assert (rdbk == 32'd11121) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                710   :   assert (rdbk == 32'd251) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                711   :   assert (rdbk == 32'd1672) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                712   :   assert (rdbk == 32'd3095) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                713   :   assert (rdbk == 32'd4520) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                714   :   assert (rdbk == 32'd5947) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                715   :   assert (rdbk == 32'd7376) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                716   :   assert (rdbk == 32'd8807) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                717   :   assert (rdbk == 32'd10240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                718   :   assert (rdbk == 32'd11675) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                719   :   assert (rdbk == 32'd823) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                720   :   assert (rdbk == 32'd2262) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                721   :   assert (rdbk == 32'd3703) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                722   :   assert (rdbk == 32'd5146) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                723   :   assert (rdbk == 32'd6591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                724   :   assert (rdbk == 32'd8038) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                725   :   assert (rdbk == 32'd9487) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                726   :   assert (rdbk == 32'd10938) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                727   :   assert (rdbk == 32'd102) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                728   :   assert (rdbk == 32'd1557) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                729   :   assert (rdbk == 32'd3014) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                730   :   assert (rdbk == 32'd4473) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                731   :   assert (rdbk == 32'd5934) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                732   :   assert (rdbk == 32'd7397) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                733   :   assert (rdbk == 32'd8862) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                734   :   assert (rdbk == 32'd10329) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                735   :   assert (rdbk == 32'd11798) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                736   :   assert (rdbk == 32'd980) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                737   :   assert (rdbk == 32'd2453) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                738   :   assert (rdbk == 32'd3928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                739   :   assert (rdbk == 32'd5405) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                740   :   assert (rdbk == 32'd6884) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                741   :   assert (rdbk == 32'd8365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                742   :   assert (rdbk == 32'd9848) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                743   :   assert (rdbk == 32'd11333) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                744   :   assert (rdbk == 32'd531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                745   :   assert (rdbk == 32'd2020) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                746   :   assert (rdbk == 32'd3511) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                747   :   assert (rdbk == 32'd5004) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                748   :   assert (rdbk == 32'd6499) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                749   :   assert (rdbk == 32'd7996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                750   :   assert (rdbk == 32'd9495) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                751   :   assert (rdbk == 32'd10996) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                752   :   assert (rdbk == 32'd210) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                753   :   assert (rdbk == 32'd1715) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                754   :   assert (rdbk == 32'd3222) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                755   :   assert (rdbk == 32'd4731) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                756   :   assert (rdbk == 32'd6242) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                757   :   assert (rdbk == 32'd7755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                758   :   assert (rdbk == 32'd9270) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                759   :   assert (rdbk == 32'd10787) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                760   :   assert (rdbk == 32'd17) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                761   :   assert (rdbk == 32'd1538) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                762   :   assert (rdbk == 32'd3061) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                763   :   assert (rdbk == 32'd4586) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                764   :   assert (rdbk == 32'd6113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                765   :   assert (rdbk == 32'd7642) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                766   :   assert (rdbk == 32'd9173) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                767   :   assert (rdbk == 32'd10706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                768   :   assert (rdbk == 32'd12241) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                769   :   assert (rdbk == 32'd1489) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                770   :   assert (rdbk == 32'd3028) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                771   :   assert (rdbk == 32'd4569) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                772   :   assert (rdbk == 32'd6112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                773   :   assert (rdbk == 32'd7657) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                774   :   assert (rdbk == 32'd9204) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                775   :   assert (rdbk == 32'd10753) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                776   :   assert (rdbk == 32'd15) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                777   :   assert (rdbk == 32'd1568) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                778   :   assert (rdbk == 32'd3123) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                779   :   assert (rdbk == 32'd4680) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                780   :   assert (rdbk == 32'd6239) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                781   :   assert (rdbk == 32'd7800) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                782   :   assert (rdbk == 32'd9363) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                783   :   assert (rdbk == 32'd10928) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                784   :   assert (rdbk == 32'd206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                785   :   assert (rdbk == 32'd1775) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                786   :   assert (rdbk == 32'd3346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                787   :   assert (rdbk == 32'd4919) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                788   :   assert (rdbk == 32'd6494) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                789   :   assert (rdbk == 32'd8071) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                790   :   assert (rdbk == 32'd9650) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                791   :   assert (rdbk == 32'd11231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                792   :   assert (rdbk == 32'd525) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                793   :   assert (rdbk == 32'd2110) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                794   :   assert (rdbk == 32'd3697) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                795   :   assert (rdbk == 32'd5286) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                796   :   assert (rdbk == 32'd6877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                797   :   assert (rdbk == 32'd8470) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                798   :   assert (rdbk == 32'd10065) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                799   :   assert (rdbk == 32'd11662) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                800   :   assert (rdbk == 32'd972) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                801   :   assert (rdbk == 32'd2573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                802   :   assert (rdbk == 32'd4176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                803   :   assert (rdbk == 32'd5781) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                804   :   assert (rdbk == 32'd7388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                805   :   assert (rdbk == 32'd8997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                806   :   assert (rdbk == 32'd10608) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                807   :   assert (rdbk == 32'd12221) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                808   :   assert (rdbk == 32'd1547) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                809   :   assert (rdbk == 32'd3164) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                810   :   assert (rdbk == 32'd4783) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                811   :   assert (rdbk == 32'd6404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                812   :   assert (rdbk == 32'd8027) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                813   :   assert (rdbk == 32'd9652) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                814   :   assert (rdbk == 32'd11279) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                815   :   assert (rdbk == 32'd619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                816   :   assert (rdbk == 32'd2250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                817   :   assert (rdbk == 32'd3883) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                818   :   assert (rdbk == 32'd5518) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                819   :   assert (rdbk == 32'd7155) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                820   :   assert (rdbk == 32'd8794) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                821   :   assert (rdbk == 32'd10435) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                822   :   assert (rdbk == 32'd12078) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                823   :   assert (rdbk == 32'd1434) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                824   :   assert (rdbk == 32'd3081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                825   :   assert (rdbk == 32'd4730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                826   :   assert (rdbk == 32'd6381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                827   :   assert (rdbk == 32'd8034) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                828   :   assert (rdbk == 32'd9689) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                829   :   assert (rdbk == 32'd11346) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                830   :   assert (rdbk == 32'd716) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                831   :   assert (rdbk == 32'd2377) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                832   :   assert (rdbk == 32'd4040) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                833   :   assert (rdbk == 32'd5705) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                834   :   assert (rdbk == 32'd7372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                835   :   assert (rdbk == 32'd9041) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                836   :   assert (rdbk == 32'd10712) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                837   :   assert (rdbk == 32'd96) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                838   :   assert (rdbk == 32'd1771) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                839   :   assert (rdbk == 32'd3448) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                840   :   assert (rdbk == 32'd5127) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                841   :   assert (rdbk == 32'd6808) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                842   :   assert (rdbk == 32'd8491) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                843   :   assert (rdbk == 32'd10176) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                844   :   assert (rdbk == 32'd11863) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                845   :   assert (rdbk == 32'd1263) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                846   :   assert (rdbk == 32'd2954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                847   :   assert (rdbk == 32'd4647) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                848   :   assert (rdbk == 32'd6342) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                849   :   assert (rdbk == 32'd8039) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                850   :   assert (rdbk == 32'd9738) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                851   :   assert (rdbk == 32'd11439) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                852   :   assert (rdbk == 32'd853) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                853   :   assert (rdbk == 32'd2558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                854   :   assert (rdbk == 32'd4265) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                855   :   assert (rdbk == 32'd5974) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                856   :   assert (rdbk == 32'd7685) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                857   :   assert (rdbk == 32'd9398) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                858   :   assert (rdbk == 32'd11113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                859   :   assert (rdbk == 32'd541) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                860   :   assert (rdbk == 32'd2260) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                861   :   assert (rdbk == 32'd3981) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                862   :   assert (rdbk == 32'd5704) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                863   :   assert (rdbk == 32'd7429) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                864   :   assert (rdbk == 32'd9156) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                865   :   assert (rdbk == 32'd10885) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                866   :   assert (rdbk == 32'd327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                867   :   assert (rdbk == 32'd2060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                868   :   assert (rdbk == 32'd3795) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                869   :   assert (rdbk == 32'd5532) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                870   :   assert (rdbk == 32'd7271) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                871   :   assert (rdbk == 32'd9012) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                872   :   assert (rdbk == 32'd10755) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                873   :   assert (rdbk == 32'd211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                874   :   assert (rdbk == 32'd1958) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                875   :   assert (rdbk == 32'd3707) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                876   :   assert (rdbk == 32'd5458) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                877   :   assert (rdbk == 32'd7211) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                878   :   assert (rdbk == 32'd8966) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                879   :   assert (rdbk == 32'd10723) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                880   :   assert (rdbk == 32'd193) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                881   :   assert (rdbk == 32'd1954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                882   :   assert (rdbk == 32'd3717) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                883   :   assert (rdbk == 32'd5482) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                884   :   assert (rdbk == 32'd7249) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                885   :   assert (rdbk == 32'd9018) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                886   :   assert (rdbk == 32'd10789) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                887   :   assert (rdbk == 32'd273) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                888   :   assert (rdbk == 32'd2048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                889   :   assert (rdbk == 32'd3825) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                890   :   assert (rdbk == 32'd5604) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                891   :   assert (rdbk == 32'd7385) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                892   :   assert (rdbk == 32'd9168) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                893   :   assert (rdbk == 32'd10953) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                894   :   assert (rdbk == 32'd451) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                895   :   assert (rdbk == 32'd2240) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                896   :   assert (rdbk == 32'd4031) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                897   :   assert (rdbk == 32'd5824) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                898   :   assert (rdbk == 32'd7619) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                899   :   assert (rdbk == 32'd9416) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                900   :   assert (rdbk == 32'd11215) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                901   :   assert (rdbk == 32'd727) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                902   :   assert (rdbk == 32'd2530) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                903   :   assert (rdbk == 32'd4335) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                904   :   assert (rdbk == 32'd6142) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                905   :   assert (rdbk == 32'd7951) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                906   :   assert (rdbk == 32'd9762) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                907   :   assert (rdbk == 32'd11575) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                908   :   assert (rdbk == 32'd1101) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                909   :   assert (rdbk == 32'd2918) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                910   :   assert (rdbk == 32'd4737) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                911   :   assert (rdbk == 32'd6558) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                912   :   assert (rdbk == 32'd8381) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                913   :   assert (rdbk == 32'd10206) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                914   :   assert (rdbk == 32'd12033) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                915   :   assert (rdbk == 32'd1573) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                916   :   assert (rdbk == 32'd3404) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                917   :   assert (rdbk == 32'd5237) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                918   :   assert (rdbk == 32'd7072) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                919   :   assert (rdbk == 32'd8909) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                920   :   assert (rdbk == 32'd10748) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                921   :   assert (rdbk == 32'd300) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                922   :   assert (rdbk == 32'd2143) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                923   :   assert (rdbk == 32'd3988) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                924   :   assert (rdbk == 32'd5835) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                925   :   assert (rdbk == 32'd7684) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                926   :   assert (rdbk == 32'd9535) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                927   :   assert (rdbk == 32'd11388) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                928   :   assert (rdbk == 32'd954) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                929   :   assert (rdbk == 32'd2811) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                930   :   assert (rdbk == 32'd4670) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                931   :   assert (rdbk == 32'd6531) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                932   :   assert (rdbk == 32'd8394) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                933   :   assert (rdbk == 32'd10259) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                934   :   assert (rdbk == 32'd12126) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                935   :   assert (rdbk == 32'd1706) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                936   :   assert (rdbk == 32'd3577) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                937   :   assert (rdbk == 32'd5450) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                938   :   assert (rdbk == 32'd7325) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                939   :   assert (rdbk == 32'd9202) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                940   :   assert (rdbk == 32'd11081) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                941   :   assert (rdbk == 32'd673) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                942   :   assert (rdbk == 32'd2556) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                943   :   assert (rdbk == 32'd4441) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                944   :   assert (rdbk == 32'd6328) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                945   :   assert (rdbk == 32'd8217) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                946   :   assert (rdbk == 32'd10108) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                947   :   assert (rdbk == 32'd12001) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                948   :   assert (rdbk == 32'd1607) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                949   :   assert (rdbk == 32'd3504) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                950   :   assert (rdbk == 32'd5403) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                951   :   assert (rdbk == 32'd7304) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                952   :   assert (rdbk == 32'd9207) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                953   :   assert (rdbk == 32'd11112) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                954   :   assert (rdbk == 32'd730) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                955   :   assert (rdbk == 32'd2639) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                956   :   assert (rdbk == 32'd4550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                957   :   assert (rdbk == 32'd6463) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                958   :   assert (rdbk == 32'd8378) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                959   :   assert (rdbk == 32'd10295) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                960   :   assert (rdbk == 32'd12214) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                961   :   assert (rdbk == 32'd1846) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                962   :   assert (rdbk == 32'd3769) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                963   :   assert (rdbk == 32'd5694) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                964   :   assert (rdbk == 32'd7621) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                965   :   assert (rdbk == 32'd9550) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                966   :   assert (rdbk == 32'd11481) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                967   :   assert (rdbk == 32'd1125) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                968   :   assert (rdbk == 32'd3060) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                969   :   assert (rdbk == 32'd4997) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                970   :   assert (rdbk == 32'd6936) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                971   :   assert (rdbk == 32'd8877) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                972   :   assert (rdbk == 32'd10820) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                973   :   assert (rdbk == 32'd476) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                974   :   assert (rdbk == 32'd2423) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                975   :   assert (rdbk == 32'd4372) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                976   :   assert (rdbk == 32'd6323) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                977   :   assert (rdbk == 32'd8276) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                978   :   assert (rdbk == 32'd10231) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                979   :   assert (rdbk == 32'd12188) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                980   :   assert (rdbk == 32'd1858) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                981   :   assert (rdbk == 32'd3819) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                982   :   assert (rdbk == 32'd5782) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                983   :   assert (rdbk == 32'd7747) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                984   :   assert (rdbk == 32'd9714) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                985   :   assert (rdbk == 32'd11683) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                986   :   assert (rdbk == 32'd1365) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                987   :   assert (rdbk == 32'd3338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                988   :   assert (rdbk == 32'd5313) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                989   :   assert (rdbk == 32'd7290) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                990   :   assert (rdbk == 32'd9269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                991   :   assert (rdbk == 32'd11250) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                992   :   assert (rdbk == 32'd944) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                993   :   assert (rdbk == 32'd2929) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                994   :   assert (rdbk == 32'd4916) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                995   :   assert (rdbk == 32'd6905) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                996   :   assert (rdbk == 32'd8896) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                997   :   assert (rdbk == 32'd10889) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                998   :   assert (rdbk == 32'd595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                999   :   assert (rdbk == 32'd2592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1000   :   assert (rdbk == 32'd4591) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1001   :   assert (rdbk == 32'd6592) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1002   :   assert (rdbk == 32'd8595) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1003   :   assert (rdbk == 32'd10600) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1004   :   assert (rdbk == 32'd318) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1005   :   assert (rdbk == 32'd2327) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1006   :   assert (rdbk == 32'd4338) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1007   :   assert (rdbk == 32'd6351) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1008   :   assert (rdbk == 32'd8366) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1009   :   assert (rdbk == 32'd10383) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1010   :   assert (rdbk == 32'd113) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1011   :   assert (rdbk == 32'd2134) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1012   :   assert (rdbk == 32'd4157) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1013   :   assert (rdbk == 32'd6182) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1014   :   assert (rdbk == 32'd8209) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1015   :   assert (rdbk == 32'd10238) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1016   :   assert (rdbk == 32'd12269) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1017   :   assert (rdbk == 32'd2013) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1018   :   assert (rdbk == 32'd4048) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1019   :   assert (rdbk == 32'd6085) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1020   :   assert (rdbk == 32'd8124) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1021   :   assert (rdbk == 32'd10165) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1022   :   assert (rdbk == 32'd12208) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
                1023   :   assert (rdbk == 32'd1964) else begin $fwrite(f,"Wrong Result!\n"); error_count ++; end
            endcase
        end
        
        // Measurement of Performance
        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Dilithium NTT Performance in CC : %d \n", cc_count_dilithium);
        $fwrite(f,"----------------------------------------------------------------\n");        

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Dilithium NTT (indirect) Performance in CC : %d \n", cc_count_dilithium_indirect);
        $fwrite(f,"----------------------------------------------------------------\n");  

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Dilithium INVNTT Performance in CC : %d \n", cc_count_dilithium_inv);
        $fwrite(f,"----------------------------------------------------------------\n");  

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Dilithium INVNTT (indirect) Performance in CC : %d \n", cc_count_dilithium_inv_indirect);
        $fwrite(f,"----------------------------------------------------------------\n"); 
        
        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Dilithium Multiplication Performance in CC : %d \n", cc_count_dilithium_pointwise_mul);
        $fwrite(f,"----------------------------------------------------------------\n");  

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Kyber NTT Performance in CC : %d \n", cc_count_kyber);
        $fwrite(f,"----------------------------------------------------------------\n");         

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Kyber INVNTT Performance in CC : %d \n", cc_count_kyber_inv);
        $fwrite(f,"----------------------------------------------------------------\n");      

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Kyber NTT (indirect)  Performance in CC : %d \n", cc_count_kyber_indirect);
        $fwrite(f,"----------------------------------------------------------------\n");  

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Kyber INVNTT (indirect) Performance in CC : %d \n", cc_count_kyber_inv_indirect);
        $fwrite(f,"----------------------------------------------------------------\n"); 

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Kyber Multiplication Performance in CC : %d \n", cc_count_kyber_base_mul);
        $fwrite(f,"----------------------------------------------------------------\n");  
 
        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-512 NTT (indirect) Performance in CC : %d \n", cc_count_falcon512_indirect);
        $fwrite(f,"----------------------------------------------------------------\n");   

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-512 INVNTT (indirect) Performance in CC : %d \n", cc_count_falcon512_inv_indirect);
        $fwrite(f,"----------------------------------------------------------------\n"); 

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-512 Multiplication Performance in CC : %d \n", cc_count_falcon512_pointwise_mul);
        $fwrite(f,"----------------------------------------------------------------\n");  

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-1024 NTT (indirect) Performance in CC : %d \n", cc_count_falcon1024_indirect);
        $fwrite(f,"----------------------------------------------------------------\n");   

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-1024 INVNTT (indirect) Performance in CC : %d \n", cc_count_falcon1024_inv_indirect);
        $fwrite(f,"----------------------------------------------------------------\n"); 

        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"FALCON-1024 Multiplication Performance in CC : %d \n", cc_count_falcon1024_pointwise_mul);
        $fwrite(f,"----------------------------------------------------------------\n");  
        
        $fwrite(f,"----------------------------------------------------------------\n");           
        $fwrite(f,"Errors: %d \n",error_count);
        $fwrite(f,"----------------------------------------------------------------\n");  
        
         
        $fclose(f);
    end
 
    assign ram_cfg_i.ram_cfg.cfg_en = 1'b0;
    assign ram_cfg_i.ram_cfg.cfg = 4'b0;   
    assign ram_cfg_i.rf_cfg.cfg_en = 1'b0;
    assign ram_cfg_i.rf_cfg.cfg = 4'b0; 
       
    assign alert_rx_i[0].ack_n  = 1'b1;
    assign alert_rx_i[0].ack_p  = 1'b0;
    assign alert_rx_i[0].ping_n = 1'b1;
    assign alert_rx_i[0].ping_p = 1'b0;
    assign alert_rx_i[1].ack_n  = 1'b1;
    assign alert_rx_i[1].ack_p  = 1'b0;
    assign alert_rx_i[1].ping_n = 1'b1;
    assign alert_rx_i[1].ping_p = 1'b0;
  
   // Generate integrity signals for bus
  // to otbn
  assign tl_i_d.a_param = 3'b0;

  assign tl_i_d.d_ready = 1'b1;
  
  tlul_cmd_intg_gen u_tlul_cmd_intg_gen (
      .tl_i(tl_i_d),
      .tl_o(tl_i_q)
  );

  // Check integrity of transmission from
  // otbn
  tlul_rsp_intg_chk u_tlul_rsp_intg_chk (
      .tl_i (tl_o),
      .err_o(err_tl)
  );
   
endmodule
